library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use STD.textio.all;
use work.debugtools.all;
use work.cputypes.all;

entity test_hyperram16 is
end entity;

architecture foo of test_hyperram16 is

  signal cpuclock : std_logic := '1';
  signal pixelclock : std_logic := '1';
  signal clock163 : std_logic := '1';
  signal clock325 : std_logic := '1';

  signal expansionram_current_cache_line_next_toggle : std_logic := '0';
  signal expansionram_read : std_logic;
  signal expansionram_write : std_logic := '0';
  signal expansionram_rdata : unsigned(15 downto 0);
  signal expansionram_wdata : unsigned(15 downto 0) := x"4242";
  signal expansionram_address : unsigned(26 downto 0) := "000000100100011010001010111";
  signal expansionram_data_ready_strobe : std_logic;
  signal expansionram_busy : std_logic;
  signal current_cache_line : cache_row_t := (others => (others => '0'));
  signal current_cache_line_address : unsigned(26 downto 3) := (others => '0');
  signal current_cache_line_valid : std_logic := '0';

  signal cycles : integer := 0;  
  
  signal slow_prefetched_address : unsigned(26 downto 0);
  signal slow_prefetched_data : unsigned(7 downto 0);
  signal slow_prefetched_request_toggle : std_logic := '0';
  
  signal hr_d : unsigned(7 downto 0) := (others => '0');
  signal hr_rwds : std_logic := '0';
  signal hr_reset : std_logic := '1';
  signal hr_clk_n : std_logic := '0';
  signal hr_clk_p : std_logic := '0';
  signal hr_cs0 : std_logic := '0';

  signal hr2_d : unsigned(7 downto 0) := (others => '0');
  signal hr2_rwds : std_logic := '0';
  signal hr2_reset : std_logic := '1';
  signal hr2_clk_n : std_logic := '0';
  signal hr2_clk_p : std_logic := '0';
  signal hr2_cs0 : std_logic := '0';
  
  type mem_transaction_t is record
    address : unsigned(27 downto 0);
    write_p : std_logic;
    value : unsigned(15 downto 0);     -- either to write, or expected to read
  end record mem_transaction_t;

  type mem_job_list_t is array(0 to 2047) of mem_transaction_t;

  signal start_time : integer := 0;
  signal current_time : integer := 0;
  signal dispatch_time : integer := 0;
  
  signal mem_jobs : mem_job_list_t := (
    -- Simple write and then read immediately
    (address => x"8801000", write_p => '1', value => x"1984"),
    (address => x"8801000", write_p => '0', value => x"1984"),

    -- Try to reproduce the read-strobe bug
    (address => x"8801000", write_p => '1', value => x"1984"),
    (address => x"8801000", write_p => '1', value => x"1984"),

    (address => x"8802000", write_p => '1', value => x"1241"),
    (address => x"8802002", write_p => '1', value => x"2342"),
    (address => x"8802004", write_p => '1', value => x"3433"),
    (address => x"8802006", write_p => '1', value => x"4534"),
    (address => x"8802008", write_p => '1', value => x"5625"),
    (address => x"8802010", write_p => '1', value => x"6726"),
    (address => x"8802012", write_p => '1', value => x"7817"),
    (address => x"8802014", write_p => '1', value => x"8918"),
    
    (address => x"8802000", write_p => '0', value => x"1241"),
    (address => x"8802002", write_p => '0', value => x"2342"),
    (address => x"8802004", write_p => '0', value => x"3433"),
    (address => x"8802006", write_p => '0', value => x"4534"),
    (address => x"8802008", write_p => '0', value => x"5625"),
    (address => x"8802010", write_p => '0', value => x"6726"),
    (address => x"8802012", write_p => '0', value => x"7817"),
    (address => x"8802014", write_p => '0', value => x"8918"),
    
    -- Issue #280, let's write then read a few pages of data, and see if we get
    -- the wrong results at the start of each page.
    -- sy2002 wrote at word $333333 onwards = real address $8666666 for us
    (address => x"8000000", write_p => '1', value => x"1234"),
    (address => x"8000000", write_p => '1', value => x"5678"),
    (address => x"8000000", write_p => '1', value => x"9abc"),
    (address => x"8666666", write_p => '1', value => x"0000"),
    (address => x"8666668", write_p => '1', value => x"0001"),
    (address => x"866666a", write_p => '1', value => x"0002"),
    (address => x"866666c", write_p => '1', value => x"0003"),
    (address => x"866666e", write_p => '1', value => x"0004"),
    (address => x"8666670", write_p => '1', value => x"0005"),
    (address => x"8666672", write_p => '1', value => x"0006"),
    (address => x"8666674", write_p => '1', value => x"0007"),
    (address => x"8666676", write_p => '1', value => x"0008"),
    (address => x"8666678", write_p => '1', value => x"0009"),
    (address => x"866667a", write_p => '1', value => x"000a"),
    (address => x"866667c", write_p => '1', value => x"000b"),
    (address => x"866667e", write_p => '1', value => x"000c"),
    (address => x"8666680", write_p => '1', value => x"000d"),
    (address => x"8666682", write_p => '1', value => x"000e"),
    (address => x"8666684", write_p => '1', value => x"000f"),
    (address => x"8666686", write_p => '1', value => x"0010"),
    (address => x"8666688", write_p => '1', value => x"0011"),
    (address => x"866668a", write_p => '1', value => x"0012"),
    (address => x"866668c", write_p => '1', value => x"0013"),
    (address => x"866668e", write_p => '1', value => x"0014"),
    (address => x"8666690", write_p => '1', value => x"0015"),
    (address => x"8666692", write_p => '1', value => x"0016"),
    (address => x"8666694", write_p => '1', value => x"0017"),
    (address => x"8666696", write_p => '1', value => x"0018"),
    (address => x"8666698", write_p => '1', value => x"0019"),
    (address => x"866669a", write_p => '1', value => x"001a"),
    (address => x"866669c", write_p => '1', value => x"001b"),
    (address => x"866669e", write_p => '1', value => x"001c"),
    (address => x"86666a0", write_p => '1', value => x"001d"),
    (address => x"86666a2", write_p => '1', value => x"001e"),
    (address => x"86666a4", write_p => '1', value => x"001f"),
    (address => x"86666a6", write_p => '1', value => x"0020"),
    (address => x"86666a8", write_p => '1', value => x"0021"),
    (address => x"86666aa", write_p => '1', value => x"0022"),
    (address => x"86666ac", write_p => '1', value => x"0023"),
    (address => x"86666ae", write_p => '1', value => x"0024"),
    (address => x"86666b0", write_p => '1', value => x"0025"),
    (address => x"86666b2", write_p => '1', value => x"0026"),
    (address => x"86666b4", write_p => '1', value => x"0027"),
    (address => x"86666b6", write_p => '1', value => x"0028"),
    (address => x"86666b8", write_p => '1', value => x"0029"),
    (address => x"86666ba", write_p => '1', value => x"002a"),
    (address => x"86666bc", write_p => '1', value => x"002b"),
    (address => x"86666be", write_p => '1', value => x"002c"),
    (address => x"86666c0", write_p => '1', value => x"002d"),
    (address => x"86666c2", write_p => '1', value => x"002e"),
    (address => x"86666c4", write_p => '1', value => x"002f"),
    (address => x"86666c6", write_p => '1', value => x"0030"),
    (address => x"86666c8", write_p => '1', value => x"0031"),
    (address => x"86666ca", write_p => '1', value => x"0032"),
    (address => x"86666cc", write_p => '1', value => x"0033"),
    (address => x"86666ce", write_p => '1', value => x"0034"),
    (address => x"86666d0", write_p => '1', value => x"0035"),
    (address => x"86666d2", write_p => '1', value => x"0036"),
    (address => x"86666d4", write_p => '1', value => x"0037"),
    (address => x"86666d6", write_p => '1', value => x"0038"),
    (address => x"86666d8", write_p => '1', value => x"0039"),
    (address => x"86666da", write_p => '1', value => x"003a"),
    (address => x"86666dc", write_p => '1', value => x"003b"),
    (address => x"86666de", write_p => '1', value => x"003c"),
    (address => x"86666e0", write_p => '1', value => x"003d"),
    (address => x"86666e2", write_p => '1', value => x"003e"),
    (address => x"86666e4", write_p => '1', value => x"003f"),
    (address => x"86666e6", write_p => '1', value => x"0040"),
    (address => x"86666e8", write_p => '1', value => x"0041"),
    (address => x"86666ea", write_p => '1', value => x"0042"),
    (address => x"86666ec", write_p => '1', value => x"0043"),
    (address => x"86666ee", write_p => '1', value => x"0044"),
    (address => x"86666f0", write_p => '1', value => x"0045"),
    (address => x"86666f2", write_p => '1', value => x"0046"),
    (address => x"86666f4", write_p => '1', value => x"0047"),
    (address => x"86666f6", write_p => '1', value => x"0048"),
    (address => x"86666f8", write_p => '1', value => x"0049"),
    (address => x"86666fa", write_p => '1', value => x"004a"),
    (address => x"86666fc", write_p => '1', value => x"004b"),
    (address => x"86666fe", write_p => '1', value => x"004c"),
    (address => x"8666700", write_p => '1', value => x"004d"),
    (address => x"8666702", write_p => '1', value => x"004e"),
    (address => x"8666704", write_p => '1', value => x"004f"),
    (address => x"8666706", write_p => '1', value => x"0050"),
    (address => x"8666708", write_p => '1', value => x"0051"),
    (address => x"866670a", write_p => '1', value => x"0052"),
    (address => x"866670c", write_p => '1', value => x"0053"),
    (address => x"866670e", write_p => '1', value => x"0054"),
    (address => x"8666710", write_p => '1', value => x"0055"),
    (address => x"8666712", write_p => '1', value => x"0056"),
    (address => x"8666714", write_p => '1', value => x"0057"),
    (address => x"8666716", write_p => '1', value => x"0058"),
    (address => x"8666718", write_p => '1', value => x"0059"),
    (address => x"866671a", write_p => '1', value => x"005a"),
    (address => x"866671c", write_p => '1', value => x"005b"),
    (address => x"866671e", write_p => '1', value => x"005c"),
    (address => x"8666720", write_p => '1', value => x"005d"),
    (address => x"8666722", write_p => '1', value => x"005e"),
    (address => x"8666724", write_p => '1', value => x"005f"),
    (address => x"8666726", write_p => '1', value => x"0060"),
    (address => x"8666728", write_p => '1', value => x"0061"),
    (address => x"866672a", write_p => '1', value => x"0062"),
    (address => x"866672c", write_p => '1', value => x"0063"),
    (address => x"866672e", write_p => '1', value => x"0064"),
    (address => x"8666730", write_p => '1', value => x"0065"),
    (address => x"8666732", write_p => '1', value => x"0066"),
    (address => x"8666734", write_p => '1', value => x"0067"),
    (address => x"8666736", write_p => '1', value => x"0068"),
    (address => x"8666738", write_p => '1', value => x"0069"),
    (address => x"866673a", write_p => '1', value => x"006a"),
    (address => x"866673c", write_p => '1', value => x"006b"),
    (address => x"866673e", write_p => '1', value => x"006c"),
    (address => x"8666740", write_p => '1', value => x"006d"),
    (address => x"8666742", write_p => '1', value => x"006e"),
    (address => x"8666744", write_p => '1', value => x"006f"),
    (address => x"8666746", write_p => '1', value => x"0070"),
    (address => x"8666748", write_p => '1', value => x"0071"),
    (address => x"866674a", write_p => '1', value => x"0072"),
    (address => x"866674c", write_p => '1', value => x"0073"),
    (address => x"866674e", write_p => '1', value => x"0074"),
    (address => x"8666750", write_p => '1', value => x"0075"),
    (address => x"8666752", write_p => '1', value => x"0076"),
    (address => x"8666754", write_p => '1', value => x"0077"),
    (address => x"8666756", write_p => '1', value => x"0078"),
    (address => x"8666758", write_p => '1', value => x"0079"),
    (address => x"866675a", write_p => '1', value => x"007a"),
    (address => x"866675c", write_p => '1', value => x"007b"),
    (address => x"866675e", write_p => '1', value => x"007c"),
    (address => x"8666760", write_p => '1', value => x"007d"),
    (address => x"8666762", write_p => '1', value => x"007e"),
    (address => x"8666764", write_p => '1', value => x"007f"),
    (address => x"8666766", write_p => '1', value => x"0080"),
    (address => x"8666768", write_p => '1', value => x"0081"),
    (address => x"866676a", write_p => '1', value => x"0082"),
    (address => x"866676c", write_p => '1', value => x"0083"),
    (address => x"866676e", write_p => '1', value => x"0084"),
    (address => x"8666770", write_p => '1', value => x"0085"),
    (address => x"8666772", write_p => '1', value => x"0086"),
    (address => x"8666774", write_p => '1', value => x"0087"),
    (address => x"8666776", write_p => '1', value => x"0088"),
    (address => x"8666778", write_p => '1', value => x"0089"),
    (address => x"866677a", write_p => '1', value => x"008a"),
    (address => x"866677c", write_p => '1', value => x"008b"),
    (address => x"866677e", write_p => '1', value => x"008c"),
    (address => x"8666780", write_p => '1', value => x"008d"),
    (address => x"8666782", write_p => '1', value => x"008e"),
    (address => x"8666784", write_p => '1', value => x"008f"),
    (address => x"8666786", write_p => '1', value => x"0090"),
    (address => x"8666788", write_p => '1', value => x"0091"),
    (address => x"866678a", write_p => '1', value => x"0092"),
    (address => x"866678c", write_p => '1', value => x"0093"),
    (address => x"866678e", write_p => '1', value => x"0094"),
    (address => x"8666790", write_p => '1', value => x"0095"),
    (address => x"8666792", write_p => '1', value => x"0096"),
    (address => x"8666794", write_p => '1', value => x"0097"),
    (address => x"8666796", write_p => '1', value => x"0098"),
    (address => x"8666798", write_p => '1', value => x"0099"),
    (address => x"866679a", write_p => '1', value => x"009a"),
    (address => x"866679c", write_p => '1', value => x"009b"),
    (address => x"866679e", write_p => '1', value => x"009c"),
    (address => x"86667a0", write_p => '1', value => x"009d"),
    (address => x"86667a2", write_p => '1', value => x"009e"),
    (address => x"86667a4", write_p => '1', value => x"009f"),
    (address => x"86667a6", write_p => '1', value => x"00a0"),
    (address => x"86667a8", write_p => '1', value => x"00a1"),
    (address => x"86667aa", write_p => '1', value => x"00a2"),
    (address => x"86667ac", write_p => '1', value => x"00a3"),
    (address => x"86667ae", write_p => '1', value => x"00a4"),
    (address => x"86667b0", write_p => '1', value => x"00a5"),
    (address => x"86667b2", write_p => '1', value => x"00a6"),
    (address => x"86667b4", write_p => '1', value => x"00a7"),
    (address => x"86667b6", write_p => '1', value => x"00a8"),
    (address => x"86667b8", write_p => '1', value => x"00a9"),
    (address => x"86667ba", write_p => '1', value => x"00aa"),
    (address => x"86667bc", write_p => '1', value => x"00ab"),
    (address => x"86667be", write_p => '1', value => x"00ac"),
    (address => x"86667c0", write_p => '1', value => x"00ad"),
    (address => x"86667c2", write_p => '1', value => x"00ae"),
    (address => x"86667c4", write_p => '1', value => x"00af"),
    (address => x"86667c6", write_p => '1', value => x"00b0"),
    (address => x"86667c8", write_p => '1', value => x"00b1"),
    (address => x"86667ca", write_p => '1', value => x"00b2"),
    (address => x"86667cc", write_p => '1', value => x"00b3"),
    (address => x"86667ce", write_p => '1', value => x"00b4"),
    (address => x"86667d0", write_p => '1', value => x"00b5"),
    (address => x"86667d2", write_p => '1', value => x"00b6"),
    (address => x"86667d4", write_p => '1', value => x"00b7"),
    (address => x"86667d6", write_p => '1', value => x"00b8"),
    (address => x"86667d8", write_p => '1', value => x"00b9"),
    (address => x"86667da", write_p => '1', value => x"00ba"),
    (address => x"86667dc", write_p => '1', value => x"00bb"),
    (address => x"86667de", write_p => '1', value => x"00bc"),
    (address => x"86667e0", write_p => '1', value => x"00bd"),
    (address => x"86667e2", write_p => '1', value => x"00be"),
    (address => x"86667e4", write_p => '1', value => x"00bf"),
    (address => x"86667e6", write_p => '1', value => x"00c0"),
    (address => x"86667e8", write_p => '1', value => x"00c1"),
    (address => x"86667ea", write_p => '1', value => x"00c2"),
    (address => x"86667ec", write_p => '1', value => x"00c3"),
    (address => x"86667ee", write_p => '1', value => x"00c4"),
    (address => x"86667f0", write_p => '1', value => x"00c5"),
    (address => x"86667f2", write_p => '1', value => x"00c6"),
    (address => x"86667f4", write_p => '1', value => x"00c7"),
    (address => x"86667f6", write_p => '1', value => x"00c8"),
    (address => x"86667f8", write_p => '1', value => x"00c9"),
    (address => x"86667fa", write_p => '1', value => x"00ca"),
    (address => x"86667fc", write_p => '1', value => x"00cb"),
    (address => x"86667fe", write_p => '1', value => x"00cc"),
    (address => x"8666800", write_p => '1', value => x"00cd"),
    (address => x"8666802", write_p => '1', value => x"00ce"),
    (address => x"8666804", write_p => '1', value => x"00cf"),
    (address => x"8666806", write_p => '1', value => x"00d0"),
    (address => x"8666808", write_p => '1', value => x"00d1"),
    (address => x"866680a", write_p => '1', value => x"00d2"),
    (address => x"866680c", write_p => '1', value => x"00d3"),
    (address => x"866680e", write_p => '1', value => x"00d4"),
    (address => x"8666810", write_p => '1', value => x"00d5"),
    (address => x"8666812", write_p => '1', value => x"00d6"),
    (address => x"8666814", write_p => '1', value => x"00d7"),
    (address => x"8666816", write_p => '1', value => x"00d8"),
    (address => x"8666818", write_p => '1', value => x"00d9"),
    (address => x"866681a", write_p => '1', value => x"00da"),
    (address => x"866681c", write_p => '1', value => x"00db"),
    (address => x"866681e", write_p => '1', value => x"00dc"),
    (address => x"8666820", write_p => '1', value => x"00dd"),
    (address => x"8666822", write_p => '1', value => x"00de"),
    (address => x"8666824", write_p => '1', value => x"00df"),
    (address => x"8666826", write_p => '1', value => x"00e0"),
    (address => x"8666828", write_p => '1', value => x"00e1"),
    (address => x"866682a", write_p => '1', value => x"00e2"),
    (address => x"866682c", write_p => '1', value => x"00e3"),
    (address => x"866682e", write_p => '1', value => x"00e4"),
    (address => x"8666830", write_p => '1', value => x"00e5"),
    (address => x"8666832", write_p => '1', value => x"00e6"),
    (address => x"8666834", write_p => '1', value => x"00e7"),
    (address => x"8666836", write_p => '1', value => x"00e8"),
    (address => x"8666838", write_p => '1', value => x"00e9"),
    (address => x"866683a", write_p => '1', value => x"00ea"),
    (address => x"866683c", write_p => '1', value => x"00eb"),
    (address => x"866683e", write_p => '1', value => x"00ec"),
    (address => x"8666840", write_p => '1', value => x"00ed"),
    (address => x"8666842", write_p => '1', value => x"00ee"),
    (address => x"8666844", write_p => '1', value => x"00ef"),
    (address => x"8666846", write_p => '1', value => x"00f0"),
    (address => x"8666848", write_p => '1', value => x"00f1"),
    (address => x"866684a", write_p => '1', value => x"00f2"),
    (address => x"866684c", write_p => '1', value => x"00f3"),
    (address => x"866684e", write_p => '1', value => x"00f4"),
    (address => x"8666850", write_p => '1', value => x"00f5"),
    (address => x"8666852", write_p => '1', value => x"00f6"),
    (address => x"8666854", write_p => '1', value => x"00f7"),
    (address => x"8666856", write_p => '1', value => x"00f8"),
    (address => x"8666858", write_p => '1', value => x"00f9"),
    (address => x"866685a", write_p => '1', value => x"00fa"),
    (address => x"866685c", write_p => '1', value => x"00fb"),
    (address => x"866685e", write_p => '1', value => x"00fc"),
    (address => x"8666860", write_p => '1', value => x"00fd"),
    (address => x"8666862", write_p => '1', value => x"00fe"),
    (address => x"8666864", write_p => '1', value => x"00ff"),
    (address => x"8666866", write_p => '1', value => x"0100"),
    (address => x"8666868", write_p => '1', value => x"0101"),
    (address => x"866686a", write_p => '1', value => x"0102"),
    (address => x"866686c", write_p => '1', value => x"0103"),
    (address => x"866686e", write_p => '1', value => x"0104"),
    (address => x"8666870", write_p => '1', value => x"0105"),
    (address => x"8666872", write_p => '1', value => x"0106"),
    (address => x"8666874", write_p => '1', value => x"0107"),
    (address => x"8666876", write_p => '1', value => x"0108"),
    (address => x"8666878", write_p => '1', value => x"0109"),
    (address => x"866687a", write_p => '1', value => x"010a"),
    (address => x"866687c", write_p => '1', value => x"010b"),
    (address => x"866687e", write_p => '1', value => x"010c"),
    (address => x"8666880", write_p => '1', value => x"010d"),
    (address => x"8666882", write_p => '1', value => x"010e"),
    (address => x"8666884", write_p => '1', value => x"010f"),
    (address => x"8666886", write_p => '1', value => x"0110"),
    (address => x"8666888", write_p => '1', value => x"0111"),
    (address => x"866688a", write_p => '1', value => x"0112"),
    (address => x"866688c", write_p => '1', value => x"0113"),
    (address => x"866688e", write_p => '1', value => x"0114"),
    (address => x"8666890", write_p => '1', value => x"0115"),
    (address => x"8666892", write_p => '1', value => x"0116"),
    (address => x"8666894", write_p => '1', value => x"0117"),
    (address => x"8666896", write_p => '1', value => x"0118"),
    (address => x"8666898", write_p => '1', value => x"0119"),
    (address => x"866689a", write_p => '1', value => x"011a"),
    (address => x"866689c", write_p => '1', value => x"011b"),
    (address => x"866689e", write_p => '1', value => x"011c"),
    (address => x"86668a0", write_p => '1', value => x"011d"),
    (address => x"86668a2", write_p => '1', value => x"011e"),
    (address => x"86668a4", write_p => '1', value => x"011f"),
    (address => x"86668a6", write_p => '1', value => x"0120"),
    (address => x"86668a8", write_p => '1', value => x"0121"),
    (address => x"86668aa", write_p => '1', value => x"0122"),
    (address => x"86668ac", write_p => '1', value => x"0123"),
    (address => x"86668ae", write_p => '1', value => x"0124"),
    (address => x"86668b0", write_p => '1', value => x"0125"),
    (address => x"86668b2", write_p => '1', value => x"0126"),
    (address => x"86668b4", write_p => '1', value => x"0127"),
    (address => x"86668b6", write_p => '1', value => x"0128"),
    (address => x"86668b8", write_p => '1', value => x"0129"),
    (address => x"86668ba", write_p => '1', value => x"012a"),
    (address => x"86668bc", write_p => '1', value => x"012b"),
    (address => x"86668be", write_p => '1', value => x"012c"),
    (address => x"86668c0", write_p => '1', value => x"012d"),
    (address => x"86668c2", write_p => '1', value => x"012e"),
    (address => x"86668c4", write_p => '1', value => x"012f"),
    (address => x"86668c6", write_p => '1', value => x"0130"),
    (address => x"86668c8", write_p => '1', value => x"0131"),
    (address => x"86668ca", write_p => '1', value => x"0132"),
    (address => x"86668cc", write_p => '1', value => x"0133"),
    (address => x"86668ce", write_p => '1', value => x"0134"),
    (address => x"86668d0", write_p => '1', value => x"0135"),
    (address => x"86668d2", write_p => '1', value => x"0136"),
    (address => x"86668d4", write_p => '1', value => x"0137"),
    (address => x"86668d6", write_p => '1', value => x"0138"),
    (address => x"86668d8", write_p => '1', value => x"0139"),
    (address => x"86668da", write_p => '1', value => x"013a"),
    (address => x"86668dc", write_p => '1', value => x"013b"),
    (address => x"86668de", write_p => '1', value => x"013c"),
    (address => x"86668e0", write_p => '1', value => x"013d"),
    (address => x"86668e2", write_p => '1', value => x"013e"),
    (address => x"86668e4", write_p => '1', value => x"013f"),
    (address => x"86668e6", write_p => '1', value => x"0140"),
    (address => x"86668e8", write_p => '1', value => x"0141"),
    (address => x"86668ea", write_p => '1', value => x"0142"),
    (address => x"86668ec", write_p => '1', value => x"0143"),
    (address => x"86668ee", write_p => '1', value => x"0144"),
    (address => x"86668f0", write_p => '1', value => x"0145"),
    (address => x"86668f2", write_p => '1', value => x"0146"),
    (address => x"86668f4", write_p => '1', value => x"0147"),
    (address => x"86668f6", write_p => '1', value => x"0148"),
    (address => x"86668f8", write_p => '1', value => x"0149"),
    (address => x"86668fa", write_p => '1', value => x"014a"),
    (address => x"86668fc", write_p => '1', value => x"014b"),
    (address => x"86668fe", write_p => '1', value => x"014c"),
    (address => x"8666900", write_p => '1', value => x"014d"),
    (address => x"8666902", write_p => '1', value => x"014e"),
    (address => x"8666904", write_p => '1', value => x"014f"),
    (address => x"8666906", write_p => '1', value => x"0150"),
    (address => x"8666908", write_p => '1', value => x"0151"),
    (address => x"866690a", write_p => '1', value => x"0152"),
    (address => x"866690c", write_p => '1', value => x"0153"),
    (address => x"866690e", write_p => '1', value => x"0154"),
    (address => x"8666910", write_p => '1', value => x"0155"),
    (address => x"8666912", write_p => '1', value => x"0156"),
    (address => x"8666914", write_p => '1', value => x"0157"),
    (address => x"8666916", write_p => '1', value => x"0158"),
    (address => x"8666918", write_p => '1', value => x"0159"),
    (address => x"866691a", write_p => '1', value => x"015a"),
    (address => x"866691c", write_p => '1', value => x"015b"),
    (address => x"866691e", write_p => '1', value => x"015c"),
    (address => x"8666920", write_p => '1', value => x"015d"),
    (address => x"8666922", write_p => '1', value => x"015e"),
    (address => x"8666924", write_p => '1', value => x"015f"),
    (address => x"8666926", write_p => '1', value => x"0160"),
    (address => x"8666928", write_p => '1', value => x"0161"),
    (address => x"866692a", write_p => '1', value => x"0162"),
    (address => x"866692c", write_p => '1', value => x"0163"),
    (address => x"866692e", write_p => '1', value => x"0164"),
    (address => x"8666930", write_p => '1', value => x"0165"),
    (address => x"8666932", write_p => '1', value => x"0166"),
    (address => x"8666934", write_p => '1', value => x"0167"),
    (address => x"8666936", write_p => '1', value => x"0168"),
    (address => x"8666938", write_p => '1', value => x"0169"),
    (address => x"866693a", write_p => '1', value => x"016a"),
    (address => x"866693c", write_p => '1', value => x"016b"),
    (address => x"866693e", write_p => '1', value => x"016c"),
    (address => x"8666940", write_p => '1', value => x"016d"),
    (address => x"8666942", write_p => '1', value => x"016e"),
    (address => x"8666944", write_p => '1', value => x"016f"),
    (address => x"8666946", write_p => '1', value => x"0170"),
    (address => x"8666948", write_p => '1', value => x"0171"),
    (address => x"866694a", write_p => '1', value => x"0172"),
    (address => x"866694c", write_p => '1', value => x"0173"),
    (address => x"866694e", write_p => '1', value => x"0174"),
    (address => x"8666950", write_p => '1', value => x"0175"),
    (address => x"8666952", write_p => '1', value => x"0176"),
    (address => x"8666954", write_p => '1', value => x"0177"),
    (address => x"8666956", write_p => '1', value => x"0178"),
    (address => x"8666958", write_p => '1', value => x"0179"),
    (address => x"866695a", write_p => '1', value => x"017a"),
    (address => x"866695c", write_p => '1', value => x"017b"),
    (address => x"866695e", write_p => '1', value => x"017c"),
    (address => x"8666960", write_p => '1', value => x"017d"),
    (address => x"8666962", write_p => '1', value => x"017e"),
    (address => x"8666964", write_p => '1', value => x"017f"),
    (address => x"8666966", write_p => '1', value => x"0180"),
    (address => x"8666968", write_p => '1', value => x"0181"),
    (address => x"866696a", write_p => '1', value => x"0182"),
    (address => x"866696c", write_p => '1', value => x"0183"),
    (address => x"866696e", write_p => '1', value => x"0184"),
    (address => x"8666970", write_p => '1', value => x"0185"),
    (address => x"8666972", write_p => '1', value => x"0186"),
    (address => x"8666974", write_p => '1', value => x"0187"),
    (address => x"8666976", write_p => '1', value => x"0188"),
    (address => x"8666978", write_p => '1', value => x"0189"),
    (address => x"866697a", write_p => '1', value => x"018a"),
    (address => x"866697c", write_p => '1', value => x"018b"),
    (address => x"866697e", write_p => '1', value => x"018c"),
    (address => x"8666980", write_p => '1', value => x"018d"),
    (address => x"8666982", write_p => '1', value => x"018e"),
    (address => x"8666984", write_p => '1', value => x"018f"),
    (address => x"8666986", write_p => '1', value => x"0190"),
    (address => x"8666988", write_p => '1', value => x"0191"),
    (address => x"866698a", write_p => '1', value => x"0192"),
    (address => x"866698c", write_p => '1', value => x"0193"),
    (address => x"866698e", write_p => '1', value => x"0194"),
    (address => x"8666990", write_p => '1', value => x"0195"),
    (address => x"8666992", write_p => '1', value => x"0196"),
    (address => x"8666994", write_p => '1', value => x"0197"),
    (address => x"8666996", write_p => '1', value => x"0198"),
    (address => x"8666998", write_p => '1', value => x"0199"),
    (address => x"866699a", write_p => '1', value => x"019a"),
    (address => x"866699c", write_p => '1', value => x"019b"),
    (address => x"866699e", write_p => '1', value => x"019c"),
    (address => x"86669a0", write_p => '1', value => x"019d"),
    (address => x"86669a2", write_p => '1', value => x"019e"),
    (address => x"86669a4", write_p => '1', value => x"019f"),
    (address => x"86669a6", write_p => '1', value => x"01a0"),
    (address => x"86669a8", write_p => '1', value => x"01a1"),
    (address => x"86669aa", write_p => '1', value => x"01a2"),
    (address => x"86669ac", write_p => '1', value => x"01a3"),
    (address => x"86669ae", write_p => '1', value => x"01a4"),
    (address => x"86669b0", write_p => '1', value => x"01a5"),
    (address => x"86669b2", write_p => '1', value => x"01a6"),
    (address => x"86669b4", write_p => '1', value => x"01a7"),
    (address => x"86669b6", write_p => '1', value => x"01a8"),
    (address => x"86669b8", write_p => '1', value => x"01a9"),
    (address => x"86669ba", write_p => '1', value => x"01aa"),
    (address => x"86669bc", write_p => '1', value => x"01ab"),
    (address => x"86669be", write_p => '1', value => x"01ac"),
    (address => x"86669c0", write_p => '1', value => x"01ad"),
    (address => x"86669c2", write_p => '1', value => x"01ae"),
    (address => x"86669c4", write_p => '1', value => x"01af"),
    (address => x"86669c6", write_p => '1', value => x"01b0"),
    (address => x"86669c8", write_p => '1', value => x"01b1"),
    (address => x"86669ca", write_p => '1', value => x"01b2"),
    (address => x"86669cc", write_p => '1', value => x"01b3"),
    (address => x"86669ce", write_p => '1', value => x"01b4"),
    (address => x"86669d0", write_p => '1', value => x"01b5"),
    (address => x"86669d2", write_p => '1', value => x"01b6"),
    (address => x"86669d4", write_p => '1', value => x"01b7"),
    (address => x"86669d6", write_p => '1', value => x"01b8"),
    (address => x"86669d8", write_p => '1', value => x"01b9"),
    (address => x"86669da", write_p => '1', value => x"01ba"),
    (address => x"86669dc", write_p => '1', value => x"01bb"),
    (address => x"86669de", write_p => '1', value => x"01bc"),
    (address => x"86669e0", write_p => '1', value => x"01bd"),
    (address => x"86669e2", write_p => '1', value => x"01be"),
    (address => x"86669e4", write_p => '1', value => x"01bf"),
    (address => x"86669e6", write_p => '1', value => x"01c0"),
    (address => x"86669e8", write_p => '1', value => x"01c1"),
    (address => x"86669ea", write_p => '1', value => x"01c2"),
    (address => x"86669ec", write_p => '1', value => x"01c3"),
    (address => x"86669ee", write_p => '1', value => x"01c4"),
    (address => x"86669f0", write_p => '1', value => x"01c5"),
    (address => x"86669f2", write_p => '1', value => x"01c6"),
    (address => x"86669f4", write_p => '1', value => x"01c7"),
    (address => x"86669f6", write_p => '1', value => x"01c8"),
    (address => x"86669f8", write_p => '1', value => x"01c9"),
    (address => x"86669fa", write_p => '1', value => x"01ca"),
    (address => x"86669fc", write_p => '1', value => x"01cb"),
    (address => x"86669fe", write_p => '1', value => x"01cc"),
    (address => x"8666a00", write_p => '1', value => x"01cd"),
    (address => x"8666a02", write_p => '1', value => x"01ce"),
    (address => x"8666a04", write_p => '1', value => x"01cf"),
    (address => x"8666a06", write_p => '1', value => x"01d0"),
    (address => x"8666a08", write_p => '1', value => x"01d1"),
    (address => x"8666a0a", write_p => '1', value => x"01d2"),
    (address => x"8666a0c", write_p => '1', value => x"01d3"),
    (address => x"8666a0e", write_p => '1', value => x"01d4"),
    (address => x"8666a10", write_p => '1', value => x"01d5"),
    (address => x"8666a12", write_p => '1', value => x"01d6"),
    (address => x"8666a14", write_p => '1', value => x"01d7"),
    (address => x"8666a16", write_p => '1', value => x"01d8"),
    (address => x"8666a18", write_p => '1', value => x"01d9"),
    (address => x"8666a1a", write_p => '1', value => x"01da"),
    (address => x"8666a1c", write_p => '1', value => x"01db"),
    (address => x"8666a1e", write_p => '1', value => x"01dc"),
    (address => x"8666a20", write_p => '1', value => x"01dd"),
    (address => x"8666a22", write_p => '1', value => x"01de"),
    (address => x"8666a24", write_p => '1', value => x"01df"),
    (address => x"8666a26", write_p => '1', value => x"01e0"),
    (address => x"8666a28", write_p => '1', value => x"01e1"),
    (address => x"8666a2a", write_p => '1', value => x"01e2"),
    (address => x"8666a2c", write_p => '1', value => x"01e3"),
    (address => x"8666a2e", write_p => '1', value => x"01e4"),
    (address => x"8666a30", write_p => '1', value => x"01e5"),
    (address => x"8666a32", write_p => '1', value => x"01e6"),
    (address => x"8666a34", write_p => '1', value => x"01e7"),
    (address => x"8666a36", write_p => '1', value => x"01e8"),
    (address => x"8666a38", write_p => '1', value => x"01e9"),
    (address => x"8666a3a", write_p => '1', value => x"01ea"),
    (address => x"8666a3c", write_p => '1', value => x"01eb"),
    (address => x"8666a3e", write_p => '1', value => x"01ec"),
    (address => x"8666a40", write_p => '1', value => x"01ed"),
    (address => x"8666a42", write_p => '1', value => x"01ee"),
    (address => x"8666a44", write_p => '1', value => x"01ef"),
    (address => x"8666a46", write_p => '1', value => x"01f0"),
    (address => x"8666a48", write_p => '1', value => x"01f1"),
    (address => x"8666a4a", write_p => '1', value => x"01f2"),
    (address => x"8666a4c", write_p => '1', value => x"01f3"),
    (address => x"8666a4e", write_p => '1', value => x"01f4"),
    (address => x"8666a50", write_p => '1', value => x"01f5"),
    (address => x"8666a52", write_p => '1', value => x"01f6"),
    (address => x"8666a54", write_p => '1', value => x"01f7"),
    (address => x"8666a56", write_p => '1', value => x"01f8"),
    (address => x"8666a58", write_p => '1', value => x"01f9"),
    (address => x"8666a5a", write_p => '1', value => x"01fa"),
    (address => x"8666a5c", write_p => '1', value => x"01fb"),
    (address => x"8666a5e", write_p => '1', value => x"01fc"),
    (address => x"8666a60", write_p => '1', value => x"01fd"),
    (address => x"8666a62", write_p => '1', value => x"01fe"),
    (address => x"8666a64", write_p => '1', value => x"01ff"),
    (address => x"8666a66", write_p => '1', value => x"0200"),
    (address => x"8666a68", write_p => '1', value => x"0201"),
    (address => x"8666a6a", write_p => '1', value => x"0202"),
    (address => x"8666a6c", write_p => '1', value => x"0203"),
    (address => x"8666a6e", write_p => '1', value => x"0204"),
    (address => x"8666a70", write_p => '1', value => x"0205"),
    (address => x"8666a72", write_p => '1', value => x"0206"),
    (address => x"8666a74", write_p => '1', value => x"0207"),
    (address => x"8666a76", write_p => '1', value => x"0208"),
    (address => x"8666a78", write_p => '1', value => x"0209"),
    (address => x"8666a7a", write_p => '1', value => x"020a"),
    (address => x"8666a7c", write_p => '1', value => x"020b"),
    (address => x"8666a7e", write_p => '1', value => x"020c"),
    (address => x"8666a80", write_p => '1', value => x"020d"),
    (address => x"8666a82", write_p => '1', value => x"020e"),
    (address => x"8666a84", write_p => '1', value => x"020f"),
    (address => x"8666a86", write_p => '1', value => x"0210"),
    (address => x"8666a88", write_p => '1', value => x"0211"),
    (address => x"8666a8a", write_p => '1', value => x"0212"),
    (address => x"8666a8c", write_p => '1', value => x"0213"),
    (address => x"8666a8e", write_p => '1', value => x"0214"),
    (address => x"8666a90", write_p => '1', value => x"0215"),
    (address => x"8666a92", write_p => '1', value => x"0216"),
    (address => x"8666a94", write_p => '1', value => x"0217"),
    (address => x"8666a96", write_p => '1', value => x"0218"),
    (address => x"8666a98", write_p => '1', value => x"0219"),
    (address => x"8666a9a", write_p => '1', value => x"021a"),
    (address => x"8666a9c", write_p => '1', value => x"021b"),
    (address => x"8666a9e", write_p => '1', value => x"021c"),
    (address => x"8666aa0", write_p => '1', value => x"021d"),
    (address => x"8666aa2", write_p => '1', value => x"021e"),
    (address => x"8666aa4", write_p => '1', value => x"021f"),
    (address => x"8666aa6", write_p => '1', value => x"0220"),
    (address => x"8666aa8", write_p => '1', value => x"0221"),
    (address => x"8666aaa", write_p => '1', value => x"0222"),
    (address => x"8666aac", write_p => '1', value => x"0223"),
    (address => x"8666aae", write_p => '1', value => x"0224"),
    (address => x"8666ab0", write_p => '1', value => x"0225"),
    (address => x"8666ab2", write_p => '1', value => x"0226"),
    (address => x"8666ab4", write_p => '1', value => x"0227"),
    (address => x"8666ab6", write_p => '1', value => x"0228"),
    (address => x"8666ab8", write_p => '1', value => x"0229"),
    (address => x"8666aba", write_p => '1', value => x"022a"),
    (address => x"8666abc", write_p => '1', value => x"022b"),
    (address => x"8666abe", write_p => '1', value => x"022c"),
    (address => x"8666ac0", write_p => '1', value => x"022d"),
    (address => x"8666ac2", write_p => '1', value => x"022e"),
    (address => x"8666ac4", write_p => '1', value => x"022f"),
    (address => x"8666ac6", write_p => '1', value => x"0230"),
    (address => x"8666ac8", write_p => '1', value => x"0231"),
    (address => x"8666aca", write_p => '1', value => x"0232"),
    (address => x"8666acc", write_p => '1', value => x"0233"),
    (address => x"8666ace", write_p => '1', value => x"0234"),
    (address => x"8666ad0", write_p => '1', value => x"0235"),
    (address => x"8666ad2", write_p => '1', value => x"0236"),
    (address => x"8666ad4", write_p => '1', value => x"0237"),
    (address => x"8666ad6", write_p => '1', value => x"0238"),
    (address => x"8666ad8", write_p => '1', value => x"0239"),
    (address => x"8666ada", write_p => '1', value => x"023a"),
    (address => x"8666adc", write_p => '1', value => x"023b"),
    (address => x"8666ade", write_p => '1', value => x"023c"),
    (address => x"8666ae0", write_p => '1', value => x"023d"),
    (address => x"8666ae2", write_p => '1', value => x"023e"),
    (address => x"8666ae4", write_p => '1', value => x"023f"),
    (address => x"8666ae6", write_p => '1', value => x"0240"),
    (address => x"8666ae8", write_p => '1', value => x"0241"),
    (address => x"8666aea", write_p => '1', value => x"0242"),
    (address => x"8666aec", write_p => '1', value => x"0243"),
    (address => x"8666aee", write_p => '1', value => x"0244"),
    (address => x"8666af0", write_p => '1', value => x"0245"),
    (address => x"8666af2", write_p => '1', value => x"0246"),
    (address => x"8666af4", write_p => '1', value => x"0247"),
    (address => x"8666af6", write_p => '1', value => x"0248"),
    (address => x"8666af8", write_p => '1', value => x"0249"),
    (address => x"8666afa", write_p => '1', value => x"024a"),
    (address => x"8666afc", write_p => '1', value => x"024b"),
    (address => x"8666afe", write_p => '1', value => x"024c"),
    (address => x"8666b00", write_p => '1', value => x"024d"),
    (address => x"8666b02", write_p => '1', value => x"024e"),
    (address => x"8666b04", write_p => '1', value => x"024f"),
    (address => x"8666b06", write_p => '1', value => x"0250"),
    (address => x"8666b08", write_p => '1', value => x"0251"),
    (address => x"8666b0a", write_p => '1', value => x"0252"),
    (address => x"8666b0c", write_p => '1', value => x"0253"),
    (address => x"8666b0e", write_p => '1', value => x"0254"),
    (address => x"8666b10", write_p => '1', value => x"0255"),
    (address => x"8666b12", write_p => '1', value => x"0256"),
    (address => x"8666b14", write_p => '1', value => x"0257"),
    (address => x"8666b16", write_p => '1', value => x"0258"),
    (address => x"8666b18", write_p => '1', value => x"0259"),
    (address => x"8666b1a", write_p => '1', value => x"025a"),
    (address => x"8666b1c", write_p => '1', value => x"025b"),
    (address => x"8666b1e", write_p => '1', value => x"025c"),
    (address => x"8666b20", write_p => '1', value => x"025d"),
    (address => x"8666b22", write_p => '1', value => x"025e"),
    (address => x"8666b24", write_p => '1', value => x"025f"),
    (address => x"8666b26", write_p => '1', value => x"0260"),
    (address => x"8666b28", write_p => '1', value => x"0261"),
    (address => x"8666b2a", write_p => '1', value => x"0262"),
    (address => x"8666b2c", write_p => '1', value => x"0263"),
    (address => x"8666b2e", write_p => '1', value => x"0264"),
    (address => x"8666b30", write_p => '1', value => x"0265"),
    (address => x"8666b32", write_p => '1', value => x"0266"),
    (address => x"8666b34", write_p => '1', value => x"0267"),
    (address => x"8666b36", write_p => '1', value => x"0268"),
    (address => x"8666b38", write_p => '1', value => x"0269"),
    (address => x"8666b3a", write_p => '1', value => x"026a"),
    (address => x"8666b3c", write_p => '1', value => x"026b"),
    (address => x"8666b3e", write_p => '1', value => x"026c"),
    (address => x"8666b40", write_p => '1', value => x"026d"),
    (address => x"8666b42", write_p => '1', value => x"026e"),
    (address => x"8666b44", write_p => '1', value => x"026f"),
    (address => x"8666b46", write_p => '1', value => x"0270"),
    (address => x"8666b48", write_p => '1', value => x"0271"),
    (address => x"8666b4a", write_p => '1', value => x"0272"),
    (address => x"8666b4c", write_p => '1', value => x"0273"),
    (address => x"8666b4e", write_p => '1', value => x"0274"),
    (address => x"8666b50", write_p => '1', value => x"0275"),
    (address => x"8666b52", write_p => '1', value => x"0276"),
    (address => x"8666b54", write_p => '1', value => x"0277"),
    (address => x"8666b56", write_p => '1', value => x"0278"),
    (address => x"8666b58", write_p => '1', value => x"0279"),
    (address => x"8666b5a", write_p => '1', value => x"027a"),
    (address => x"8666b5c", write_p => '1', value => x"027b"),
    (address => x"8666b5e", write_p => '1', value => x"027c"),
    (address => x"8666b60", write_p => '1', value => x"027d"),
    (address => x"8666b62", write_p => '1', value => x"027e"),
    (address => x"8666b64", write_p => '1', value => x"027f"),
    (address => x"8666b66", write_p => '1', value => x"0280"),
    (address => x"8666b68", write_p => '1', value => x"0281"),
    (address => x"8666b6a", write_p => '1', value => x"0282"),
    (address => x"8666b6c", write_p => '1', value => x"0283"),
    (address => x"8666b6e", write_p => '1', value => x"0284"),
    (address => x"8666b70", write_p => '1', value => x"0285"),
    (address => x"8666b72", write_p => '1', value => x"0286"),
    (address => x"8666b74", write_p => '1', value => x"0287"),
    (address => x"8666b76", write_p => '1', value => x"0288"),
    (address => x"8666b78", write_p => '1', value => x"0289"),
    (address => x"8666b7a", write_p => '1', value => x"028a"),
    (address => x"8666b7c", write_p => '1', value => x"028b"),
    (address => x"8666b7e", write_p => '1', value => x"028c"),
    (address => x"8666b80", write_p => '1', value => x"028d"),
    (address => x"8666b82", write_p => '1', value => x"028e"),
    (address => x"8666b84", write_p => '1', value => x"028f"),
    (address => x"8666b86", write_p => '1', value => x"0290"),
    (address => x"8666b88", write_p => '1', value => x"0291"),
    (address => x"8666b8a", write_p => '1', value => x"0292"),
    (address => x"8666b8c", write_p => '1', value => x"0293"),
    (address => x"8666b8e", write_p => '1', value => x"0294"),
    (address => x"8666b90", write_p => '1', value => x"0295"),
    (address => x"8666b92", write_p => '1', value => x"0296"),
    (address => x"8666b94", write_p => '1', value => x"0297"),
    (address => x"8666b96", write_p => '1', value => x"0298"),
    (address => x"8666b98", write_p => '1', value => x"0299"),
    (address => x"8666b9a", write_p => '1', value => x"029a"),
    (address => x"8666b9c", write_p => '1', value => x"029b"),
    (address => x"8666b9e", write_p => '1', value => x"029c"),
    (address => x"8666ba0", write_p => '1', value => x"029d"),
    (address => x"8666ba2", write_p => '1', value => x"029e"),
    (address => x"8666ba4", write_p => '1', value => x"029f"),
    (address => x"8666ba6", write_p => '1', value => x"02a0"),
    (address => x"8666ba8", write_p => '1', value => x"02a1"),
    (address => x"8666baa", write_p => '1', value => x"02a2"),
    (address => x"8666bac", write_p => '1', value => x"02a3"),
    (address => x"8666bae", write_p => '1', value => x"02a4"),
    (address => x"8666bb0", write_p => '1', value => x"02a5"),
    (address => x"8666bb2", write_p => '1', value => x"02a6"),
    (address => x"8666bb4", write_p => '1', value => x"02a7"),
    (address => x"8666bb6", write_p => '1', value => x"02a8"),
    (address => x"8666bb8", write_p => '1', value => x"02a9"),
    (address => x"8666bba", write_p => '1', value => x"02aa"),
    (address => x"8666bbc", write_p => '1', value => x"02ab"),
    (address => x"8666bbe", write_p => '1', value => x"02ac"),
    (address => x"8666bc0", write_p => '1', value => x"02ad"),
    (address => x"8666bc2", write_p => '1', value => x"02ae"),
    (address => x"8666bc4", write_p => '1', value => x"02af"),
    (address => x"8666bc6", write_p => '1', value => x"02b0"),
    (address => x"8666bc8", write_p => '1', value => x"02b1"),
    (address => x"8666bca", write_p => '1', value => x"02b2"),
    (address => x"8666bcc", write_p => '1', value => x"02b3"),
    (address => x"8666bce", write_p => '1', value => x"02b4"),
    (address => x"8666bd0", write_p => '1', value => x"02b5"),
    (address => x"8666bd2", write_p => '1', value => x"02b6"),
    (address => x"8666bd4", write_p => '1', value => x"02b7"),
    (address => x"8666bd6", write_p => '1', value => x"02b8"),
    (address => x"8666bd8", write_p => '1', value => x"02b9"),
    (address => x"8666bda", write_p => '1', value => x"02ba"),
    (address => x"8666bdc", write_p => '1', value => x"02bb"),
    (address => x"8666bde", write_p => '1', value => x"02bc"),
    (address => x"8666be0", write_p => '1', value => x"02bd"),
    (address => x"8666be2", write_p => '1', value => x"02be"),
    (address => x"8666be4", write_p => '1', value => x"02bf"),
    (address => x"8666be6", write_p => '1', value => x"02c0"),
    (address => x"8666be8", write_p => '1', value => x"02c1"),
    (address => x"8666bea", write_p => '1', value => x"02c2"),
    (address => x"8666bec", write_p => '1', value => x"02c3"),
    (address => x"8666bee", write_p => '1', value => x"02c4"),
    (address => x"8666bf0", write_p => '1', value => x"02c5"),
    (address => x"8666bf2", write_p => '1', value => x"02c6"),
    (address => x"8666bf4", write_p => '1', value => x"02c7"),
    (address => x"8666bf6", write_p => '1', value => x"02c8"),
    (address => x"8666bf8", write_p => '1', value => x"02c9"),
    (address => x"8666bfa", write_p => '1', value => x"02ca"),
    (address => x"8666bfc", write_p => '1', value => x"02cb"),
    (address => x"8666bfe", write_p => '1', value => x"02cc"),
    (address => x"8666c00", write_p => '1', value => x"02cd"),
    (address => x"8666c02", write_p => '1', value => x"02ce"),
    (address => x"8666c04", write_p => '1', value => x"02cf"),
    (address => x"8666c06", write_p => '1', value => x"02d0"),
    (address => x"8666c08", write_p => '1', value => x"02d1"),
    (address => x"8666c0a", write_p => '1', value => x"02d2"),
    (address => x"8666c0c", write_p => '1', value => x"02d3"),
    (address => x"8666c0e", write_p => '1', value => x"02d4"),
    (address => x"8666c10", write_p => '1', value => x"02d5"),
    (address => x"8666c12", write_p => '1', value => x"02d6"),
    (address => x"8666c14", write_p => '1', value => x"02d7"),
    (address => x"8666c16", write_p => '1', value => x"02d8"),
    (address => x"8666c18", write_p => '1', value => x"02d9"),
    (address => x"8666c1a", write_p => '1', value => x"02da"),
    (address => x"8666c1c", write_p => '1', value => x"02db"),
    (address => x"8666c1e", write_p => '1', value => x"02dc"),
    (address => x"8666c20", write_p => '1', value => x"02dd"),
    (address => x"8666c22", write_p => '1', value => x"02de"),
    (address => x"8666c24", write_p => '1', value => x"02df"),
    (address => x"8666c26", write_p => '1', value => x"02e0"),
    (address => x"8666c28", write_p => '1', value => x"02e1"),
    (address => x"8666c2a", write_p => '1', value => x"02e2"),
    (address => x"8666c2c", write_p => '1', value => x"02e3"),
    (address => x"8666c2e", write_p => '1', value => x"02e4"),
    (address => x"8666c30", write_p => '1', value => x"02e5"),
    (address => x"8666c32", write_p => '1', value => x"02e6"),
    (address => x"8666c34", write_p => '1', value => x"02e7"),
    (address => x"8666c36", write_p => '1', value => x"02e8"),
    (address => x"8666c38", write_p => '1', value => x"02e9"),
    (address => x"8666c3a", write_p => '1', value => x"02ea"),
    (address => x"8666c3c", write_p => '1', value => x"02eb"),
    (address => x"8666c3e", write_p => '1', value => x"02ec"),
    (address => x"8666c40", write_p => '1', value => x"02ed"),
    (address => x"8666c42", write_p => '1', value => x"02ee"),
    (address => x"8666c44", write_p => '1', value => x"02ef"),
    (address => x"8666c46", write_p => '1', value => x"02f0"),
    (address => x"8666c48", write_p => '1', value => x"02f1"),
    (address => x"8666c4a", write_p => '1', value => x"02f2"),
    (address => x"8666c4c", write_p => '1', value => x"02f3"),
    (address => x"8666c4e", write_p => '1', value => x"02f4"),
    (address => x"8666c50", write_p => '1', value => x"02f5"),
    (address => x"8666c52", write_p => '1', value => x"02f6"),
    (address => x"8666c54", write_p => '1', value => x"02f7"),
    (address => x"8666c56", write_p => '1', value => x"02f8"),
    (address => x"8666c58", write_p => '1', value => x"02f9"),
    (address => x"8666c5a", write_p => '1', value => x"02fa"),
    (address => x"8666c5c", write_p => '1', value => x"02fb"),
    (address => x"8666c5e", write_p => '1', value => x"02fc"),
    (address => x"8666c60", write_p => '1', value => x"02fd"),
    (address => x"8666c62", write_p => '1', value => x"02fe"),
    (address => x"8666c64", write_p => '1', value => x"02ff"),
    (address => x"8666666", write_p => '0', value => x"0000"),
    (address => x"8666668", write_p => '0', value => x"0001"),
    (address => x"866666a", write_p => '0', value => x"0002"),
    (address => x"866666c", write_p => '0', value => x"0003"),
    (address => x"866666e", write_p => '0', value => x"0004"),
    (address => x"8666670", write_p => '0', value => x"0005"),
    (address => x"8666672", write_p => '0', value => x"0006"),
    (address => x"8666674", write_p => '0', value => x"0007"),
    (address => x"8666676", write_p => '0', value => x"0008"),
    (address => x"8666678", write_p => '0', value => x"0009"),
    (address => x"866667a", write_p => '0', value => x"000a"),
    (address => x"866667c", write_p => '0', value => x"000b"),
    (address => x"866667e", write_p => '0', value => x"000c"),
    (address => x"8666680", write_p => '0', value => x"000d"),
    (address => x"8666682", write_p => '0', value => x"000e"),
    (address => x"8666684", write_p => '0', value => x"000f"),
    (address => x"8666686", write_p => '0', value => x"0010"),
    (address => x"8666688", write_p => '0', value => x"0011"),
    (address => x"866668a", write_p => '0', value => x"0012"),
    (address => x"866668c", write_p => '0', value => x"0013"),
    (address => x"866668e", write_p => '0', value => x"0014"),
    (address => x"8666690", write_p => '0', value => x"0015"),
    (address => x"8666692", write_p => '0', value => x"0016"),
    (address => x"8666694", write_p => '0', value => x"0017"),
    (address => x"8666696", write_p => '0', value => x"0018"),
    (address => x"8666698", write_p => '0', value => x"0019"),
    (address => x"866669a", write_p => '0', value => x"001a"),
    (address => x"866669c", write_p => '0', value => x"001b"),
    (address => x"866669e", write_p => '0', value => x"001c"),
    (address => x"86666a0", write_p => '0', value => x"001d"),
    (address => x"86666a2", write_p => '0', value => x"001e"),
    (address => x"86666a4", write_p => '0', value => x"001f"),
    (address => x"86666a6", write_p => '0', value => x"0020"),
    (address => x"86666a8", write_p => '0', value => x"0021"),
    (address => x"86666aa", write_p => '0', value => x"0022"),
    (address => x"86666ac", write_p => '0', value => x"0023"),
    (address => x"86666ae", write_p => '0', value => x"0024"),
    (address => x"86666b0", write_p => '0', value => x"0025"),
    (address => x"86666b2", write_p => '0', value => x"0026"),
    (address => x"86666b4", write_p => '0', value => x"0027"),
    (address => x"86666b6", write_p => '0', value => x"0028"),
    (address => x"86666b8", write_p => '0', value => x"0029"),
    (address => x"86666ba", write_p => '0', value => x"002a"),
    (address => x"86666bc", write_p => '0', value => x"002b"),
    (address => x"86666be", write_p => '0', value => x"002c"),
    (address => x"86666c0", write_p => '0', value => x"002d"),
    (address => x"86666c2", write_p => '0', value => x"002e"),
    (address => x"86666c4", write_p => '0', value => x"002f"),
    (address => x"86666c6", write_p => '0', value => x"0030"),
    (address => x"86666c8", write_p => '0', value => x"0031"),
    (address => x"86666ca", write_p => '0', value => x"0032"),
    (address => x"86666cc", write_p => '0', value => x"0033"),
    (address => x"86666ce", write_p => '0', value => x"0034"),
    (address => x"86666d0", write_p => '0', value => x"0035"),
    (address => x"86666d2", write_p => '0', value => x"0036"),
    (address => x"86666d4", write_p => '0', value => x"0037"),
    (address => x"86666d6", write_p => '0', value => x"0038"),
    (address => x"86666d8", write_p => '0', value => x"0039"),
    (address => x"86666da", write_p => '0', value => x"003a"),
    (address => x"86666dc", write_p => '0', value => x"003b"),
    (address => x"86666de", write_p => '0', value => x"003c"),
    (address => x"86666e0", write_p => '0', value => x"003d"),
    (address => x"86666e2", write_p => '0', value => x"003e"),
    (address => x"86666e4", write_p => '0', value => x"003f"),
    (address => x"86666e6", write_p => '0', value => x"0040"),
    (address => x"86666e8", write_p => '0', value => x"0041"),
    (address => x"86666ea", write_p => '0', value => x"0042"),
    (address => x"86666ec", write_p => '0', value => x"0043"),
    (address => x"86666ee", write_p => '0', value => x"0044"),
    (address => x"86666f0", write_p => '0', value => x"0045"),
    (address => x"86666f2", write_p => '0', value => x"0046"),
    (address => x"86666f4", write_p => '0', value => x"0047"),
    (address => x"86666f6", write_p => '0', value => x"0048"),
    (address => x"86666f8", write_p => '0', value => x"0049"),
    (address => x"86666fa", write_p => '0', value => x"004a"),
    (address => x"86666fc", write_p => '0', value => x"004b"),
    (address => x"86666fe", write_p => '0', value => x"004c"),
    (address => x"8666700", write_p => '0', value => x"004d"),
    (address => x"8666702", write_p => '0', value => x"004e"),
    (address => x"8666704", write_p => '0', value => x"004f"),
    (address => x"8666706", write_p => '0', value => x"0050"),
    (address => x"8666708", write_p => '0', value => x"0051"),
    (address => x"866670a", write_p => '0', value => x"0052"),
    (address => x"866670c", write_p => '0', value => x"0053"),
    (address => x"866670e", write_p => '0', value => x"0054"),
    (address => x"8666710", write_p => '0', value => x"0055"),
    (address => x"8666712", write_p => '0', value => x"0056"),
    (address => x"8666714", write_p => '0', value => x"0057"),
    (address => x"8666716", write_p => '0', value => x"0058"),
    (address => x"8666718", write_p => '0', value => x"0059"),
    (address => x"866671a", write_p => '0', value => x"005a"),
    (address => x"866671c", write_p => '0', value => x"005b"),
    (address => x"866671e", write_p => '0', value => x"005c"),
    (address => x"8666720", write_p => '0', value => x"005d"),
    (address => x"8666722", write_p => '0', value => x"005e"),
    (address => x"8666724", write_p => '0', value => x"005f"),
    (address => x"8666726", write_p => '0', value => x"0060"),
    (address => x"8666728", write_p => '0', value => x"0061"),
    (address => x"866672a", write_p => '0', value => x"0062"),
    (address => x"866672c", write_p => '0', value => x"0063"),
    (address => x"866672e", write_p => '0', value => x"0064"),
    (address => x"8666730", write_p => '0', value => x"0065"),
    (address => x"8666732", write_p => '0', value => x"0066"),
    (address => x"8666734", write_p => '0', value => x"0067"),
    (address => x"8666736", write_p => '0', value => x"0068"),
    (address => x"8666738", write_p => '0', value => x"0069"),
    (address => x"866673a", write_p => '0', value => x"006a"),
    (address => x"866673c", write_p => '0', value => x"006b"),
    (address => x"866673e", write_p => '0', value => x"006c"),
    (address => x"8666740", write_p => '0', value => x"006d"),
    (address => x"8666742", write_p => '0', value => x"006e"),
    (address => x"8666744", write_p => '0', value => x"006f"),
    (address => x"8666746", write_p => '0', value => x"0070"),
    (address => x"8666748", write_p => '0', value => x"0071"),
    (address => x"866674a", write_p => '0', value => x"0072"),
    (address => x"866674c", write_p => '0', value => x"0073"),
    (address => x"866674e", write_p => '0', value => x"0074"),
    (address => x"8666750", write_p => '0', value => x"0075"),
    (address => x"8666752", write_p => '0', value => x"0076"),
    (address => x"8666754", write_p => '0', value => x"0077"),
    (address => x"8666756", write_p => '0', value => x"0078"),
    (address => x"8666758", write_p => '0', value => x"0079"),
    (address => x"866675a", write_p => '0', value => x"007a"),
    (address => x"866675c", write_p => '0', value => x"007b"),
    (address => x"866675e", write_p => '0', value => x"007c"),
    (address => x"8666760", write_p => '0', value => x"007d"),
    (address => x"8666762", write_p => '0', value => x"007e"),
    (address => x"8666764", write_p => '0', value => x"007f"),
    (address => x"8666766", write_p => '0', value => x"0080"),
    (address => x"8666768", write_p => '0', value => x"0081"),
    (address => x"866676a", write_p => '0', value => x"0082"),
    (address => x"866676c", write_p => '0', value => x"0083"),
    (address => x"866676e", write_p => '0', value => x"0084"),
    (address => x"8666770", write_p => '0', value => x"0085"),
    (address => x"8666772", write_p => '0', value => x"0086"),
    (address => x"8666774", write_p => '0', value => x"0087"),
    (address => x"8666776", write_p => '0', value => x"0088"),
    (address => x"8666778", write_p => '0', value => x"0089"),
    (address => x"866677a", write_p => '0', value => x"008a"),
    (address => x"866677c", write_p => '0', value => x"008b"),
    (address => x"866677e", write_p => '0', value => x"008c"),
    (address => x"8666780", write_p => '0', value => x"008d"),
    (address => x"8666782", write_p => '0', value => x"008e"),
    (address => x"8666784", write_p => '0', value => x"008f"),
    (address => x"8666786", write_p => '0', value => x"0090"),
    (address => x"8666788", write_p => '0', value => x"0091"),
    (address => x"866678a", write_p => '0', value => x"0092"),
    (address => x"866678c", write_p => '0', value => x"0093"),
    (address => x"866678e", write_p => '0', value => x"0094"),
    (address => x"8666790", write_p => '0', value => x"0095"),
    (address => x"8666792", write_p => '0', value => x"0096"),
    (address => x"8666794", write_p => '0', value => x"0097"),
    (address => x"8666796", write_p => '0', value => x"0098"),
    (address => x"8666798", write_p => '0', value => x"0099"),
    (address => x"866679a", write_p => '0', value => x"009a"),
    (address => x"866679c", write_p => '0', value => x"009b"),
    (address => x"866679e", write_p => '0', value => x"009c"),
    (address => x"86667a0", write_p => '0', value => x"009d"),
    (address => x"86667a2", write_p => '0', value => x"009e"),
    (address => x"86667a4", write_p => '0', value => x"009f"),
    (address => x"86667a6", write_p => '0', value => x"00a0"),
    (address => x"86667a8", write_p => '0', value => x"00a1"),
    (address => x"86667aa", write_p => '0', value => x"00a2"),
    (address => x"86667ac", write_p => '0', value => x"00a3"),
    (address => x"86667ae", write_p => '0', value => x"00a4"),
    (address => x"86667b0", write_p => '0', value => x"00a5"),
    (address => x"86667b2", write_p => '0', value => x"00a6"),
    (address => x"86667b4", write_p => '0', value => x"00a7"),
    (address => x"86667b6", write_p => '0', value => x"00a8"),
    (address => x"86667b8", write_p => '0', value => x"00a9"),
    (address => x"86667ba", write_p => '0', value => x"00aa"),
    (address => x"86667bc", write_p => '0', value => x"00ab"),
    (address => x"86667be", write_p => '0', value => x"00ac"),
    (address => x"86667c0", write_p => '0', value => x"00ad"),
    (address => x"86667c2", write_p => '0', value => x"00ae"),
    (address => x"86667c4", write_p => '0', value => x"00af"),
    (address => x"86667c6", write_p => '0', value => x"00b0"),
    (address => x"86667c8", write_p => '0', value => x"00b1"),
    (address => x"86667ca", write_p => '0', value => x"00b2"),
    (address => x"86667cc", write_p => '0', value => x"00b3"),
    (address => x"86667ce", write_p => '0', value => x"00b4"),
    (address => x"86667d0", write_p => '0', value => x"00b5"),
    (address => x"86667d2", write_p => '0', value => x"00b6"),
    (address => x"86667d4", write_p => '0', value => x"00b7"),
    (address => x"86667d6", write_p => '0', value => x"00b8"),
    (address => x"86667d8", write_p => '0', value => x"00b9"),
    (address => x"86667da", write_p => '0', value => x"00ba"),
    (address => x"86667dc", write_p => '0', value => x"00bb"),
    (address => x"86667de", write_p => '0', value => x"00bc"),
    (address => x"86667e0", write_p => '0', value => x"00bd"),
    (address => x"86667e2", write_p => '0', value => x"00be"),
    (address => x"86667e4", write_p => '0', value => x"00bf"),
    (address => x"86667e6", write_p => '0', value => x"00c0"),
    (address => x"86667e8", write_p => '0', value => x"00c1"),
    (address => x"86667ea", write_p => '0', value => x"00c2"),
    (address => x"86667ec", write_p => '0', value => x"00c3"),
    (address => x"86667ee", write_p => '0', value => x"00c4"),
    (address => x"86667f0", write_p => '0', value => x"00c5"),
    (address => x"86667f2", write_p => '0', value => x"00c6"),
    (address => x"86667f4", write_p => '0', value => x"00c7"),
    (address => x"86667f6", write_p => '0', value => x"00c8"),
    (address => x"86667f8", write_p => '0', value => x"00c9"),
    (address => x"86667fa", write_p => '0', value => x"00ca"),
    (address => x"86667fc", write_p => '0', value => x"00cb"),
    (address => x"86667fe", write_p => '0', value => x"00cc"),
    (address => x"8666800", write_p => '0', value => x"00cd"),
    (address => x"8666802", write_p => '0', value => x"00ce"),
    (address => x"8666804", write_p => '0', value => x"00cf"),
    (address => x"8666806", write_p => '0', value => x"00d0"),
    (address => x"8666808", write_p => '0', value => x"00d1"),
    (address => x"866680a", write_p => '0', value => x"00d2"),
    (address => x"866680c", write_p => '0', value => x"00d3"),
    (address => x"866680e", write_p => '0', value => x"00d4"),
    (address => x"8666810", write_p => '0', value => x"00d5"),
    (address => x"8666812", write_p => '0', value => x"00d6"),
    (address => x"8666814", write_p => '0', value => x"00d7"),
    (address => x"8666816", write_p => '0', value => x"00d8"),
    (address => x"8666818", write_p => '0', value => x"00d9"),
    (address => x"866681a", write_p => '0', value => x"00da"),
    (address => x"866681c", write_p => '0', value => x"00db"),
    (address => x"866681e", write_p => '0', value => x"00dc"),
    (address => x"8666820", write_p => '0', value => x"00dd"),
    (address => x"8666822", write_p => '0', value => x"00de"),
    (address => x"8666824", write_p => '0', value => x"00df"),
    (address => x"8666826", write_p => '0', value => x"00e0"),
    (address => x"8666828", write_p => '0', value => x"00e1"),
    (address => x"866682a", write_p => '0', value => x"00e2"),
    (address => x"866682c", write_p => '0', value => x"00e3"),
    (address => x"866682e", write_p => '0', value => x"00e4"),
    (address => x"8666830", write_p => '0', value => x"00e5"),
    (address => x"8666832", write_p => '0', value => x"00e6"),
    (address => x"8666834", write_p => '0', value => x"00e7"),
    (address => x"8666836", write_p => '0', value => x"00e8"),
    (address => x"8666838", write_p => '0', value => x"00e9"),
    (address => x"866683a", write_p => '0', value => x"00ea"),
    (address => x"866683c", write_p => '0', value => x"00eb"),
    (address => x"866683e", write_p => '0', value => x"00ec"),
    (address => x"8666840", write_p => '0', value => x"00ed"),
    (address => x"8666842", write_p => '0', value => x"00ee"),
    (address => x"8666844", write_p => '0', value => x"00ef"),
    (address => x"8666846", write_p => '0', value => x"00f0"),
    (address => x"8666848", write_p => '0', value => x"00f1"),
    (address => x"866684a", write_p => '0', value => x"00f2"),
    (address => x"866684c", write_p => '0', value => x"00f3"),
    (address => x"866684e", write_p => '0', value => x"00f4"),
    (address => x"8666850", write_p => '0', value => x"00f5"),
    (address => x"8666852", write_p => '0', value => x"00f6"),
    (address => x"8666854", write_p => '0', value => x"00f7"),
    (address => x"8666856", write_p => '0', value => x"00f8"),
    (address => x"8666858", write_p => '0', value => x"00f9"),
    (address => x"866685a", write_p => '0', value => x"00fa"),
    (address => x"866685c", write_p => '0', value => x"00fb"),
    (address => x"866685e", write_p => '0', value => x"00fc"),
    (address => x"8666860", write_p => '0', value => x"00fd"),
    (address => x"8666862", write_p => '0', value => x"00fe"),
    (address => x"8666864", write_p => '0', value => x"00ff"),
    (address => x"8666866", write_p => '0', value => x"0100"),
    (address => x"8666868", write_p => '0', value => x"0101"),
    (address => x"866686a", write_p => '0', value => x"0102"),
    (address => x"866686c", write_p => '0', value => x"0103"),
    (address => x"866686e", write_p => '0', value => x"0104"),
    (address => x"8666870", write_p => '0', value => x"0105"),
    (address => x"8666872", write_p => '0', value => x"0106"),
    (address => x"8666874", write_p => '0', value => x"0107"),
    (address => x"8666876", write_p => '0', value => x"0108"),
    (address => x"8666878", write_p => '0', value => x"0109"),
    (address => x"866687a", write_p => '0', value => x"010a"),
    (address => x"866687c", write_p => '0', value => x"010b"),
    (address => x"866687e", write_p => '0', value => x"010c"),
    (address => x"8666880", write_p => '0', value => x"010d"),
    (address => x"8666882", write_p => '0', value => x"010e"),
    (address => x"8666884", write_p => '0', value => x"010f"),
    (address => x"8666886", write_p => '0', value => x"0110"),
    (address => x"8666888", write_p => '0', value => x"0111"),
    (address => x"866688a", write_p => '0', value => x"0112"),
    (address => x"866688c", write_p => '0', value => x"0113"),
    (address => x"866688e", write_p => '0', value => x"0114"),
    (address => x"8666890", write_p => '0', value => x"0115"),
    (address => x"8666892", write_p => '0', value => x"0116"),
    (address => x"8666894", write_p => '0', value => x"0117"),
    (address => x"8666896", write_p => '0', value => x"0118"),
    (address => x"8666898", write_p => '0', value => x"0119"),
    (address => x"866689a", write_p => '0', value => x"011a"),
    (address => x"866689c", write_p => '0', value => x"011b"),
    (address => x"866689e", write_p => '0', value => x"011c"),
    (address => x"86668a0", write_p => '0', value => x"011d"),
    (address => x"86668a2", write_p => '0', value => x"011e"),
    (address => x"86668a4", write_p => '0', value => x"011f"),
    (address => x"86668a6", write_p => '0', value => x"0120"),
    (address => x"86668a8", write_p => '0', value => x"0121"),
    (address => x"86668aa", write_p => '0', value => x"0122"),
    (address => x"86668ac", write_p => '0', value => x"0123"),
    (address => x"86668ae", write_p => '0', value => x"0124"),
    (address => x"86668b0", write_p => '0', value => x"0125"),
    (address => x"86668b2", write_p => '0', value => x"0126"),
    (address => x"86668b4", write_p => '0', value => x"0127"),
    (address => x"86668b6", write_p => '0', value => x"0128"),
    (address => x"86668b8", write_p => '0', value => x"0129"),
    (address => x"86668ba", write_p => '0', value => x"012a"),
    (address => x"86668bc", write_p => '0', value => x"012b"),
    (address => x"86668be", write_p => '0', value => x"012c"),
    (address => x"86668c0", write_p => '0', value => x"012d"),
    (address => x"86668c2", write_p => '0', value => x"012e"),
    (address => x"86668c4", write_p => '0', value => x"012f"),
    (address => x"86668c6", write_p => '0', value => x"0130"),
    (address => x"86668c8", write_p => '0', value => x"0131"),
    (address => x"86668ca", write_p => '0', value => x"0132"),
    (address => x"86668cc", write_p => '0', value => x"0133"),
    (address => x"86668ce", write_p => '0', value => x"0134"),
    (address => x"86668d0", write_p => '0', value => x"0135"),
    (address => x"86668d2", write_p => '0', value => x"0136"),
    (address => x"86668d4", write_p => '0', value => x"0137"),
    (address => x"86668d6", write_p => '0', value => x"0138"),
    (address => x"86668d8", write_p => '0', value => x"0139"),
    (address => x"86668da", write_p => '0', value => x"013a"),
    (address => x"86668dc", write_p => '0', value => x"013b"),
    (address => x"86668de", write_p => '0', value => x"013c"),
    (address => x"86668e0", write_p => '0', value => x"013d"),
    (address => x"86668e2", write_p => '0', value => x"013e"),
    (address => x"86668e4", write_p => '0', value => x"013f"),
    (address => x"86668e6", write_p => '0', value => x"0140"),
    (address => x"86668e8", write_p => '0', value => x"0141"),
    (address => x"86668ea", write_p => '0', value => x"0142"),
    (address => x"86668ec", write_p => '0', value => x"0143"),
    (address => x"86668ee", write_p => '0', value => x"0144"),
    (address => x"86668f0", write_p => '0', value => x"0145"),
    (address => x"86668f2", write_p => '0', value => x"0146"),
    (address => x"86668f4", write_p => '0', value => x"0147"),
    (address => x"86668f6", write_p => '0', value => x"0148"),
    (address => x"86668f8", write_p => '0', value => x"0149"),
    (address => x"86668fa", write_p => '0', value => x"014a"),
    (address => x"86668fc", write_p => '0', value => x"014b"),
    (address => x"86668fe", write_p => '0', value => x"014c"),
    (address => x"8666900", write_p => '0', value => x"014d"),
    (address => x"8666902", write_p => '0', value => x"014e"),
    (address => x"8666904", write_p => '0', value => x"014f"),
    (address => x"8666906", write_p => '0', value => x"0150"),
    (address => x"8666908", write_p => '0', value => x"0151"),
    (address => x"866690a", write_p => '0', value => x"0152"),
    (address => x"866690c", write_p => '0', value => x"0153"),
    (address => x"866690e", write_p => '0', value => x"0154"),
    (address => x"8666910", write_p => '0', value => x"0155"),
    (address => x"8666912", write_p => '0', value => x"0156"),
    (address => x"8666914", write_p => '0', value => x"0157"),
    (address => x"8666916", write_p => '0', value => x"0158"),
    (address => x"8666918", write_p => '0', value => x"0159"),
    (address => x"866691a", write_p => '0', value => x"015a"),
    (address => x"866691c", write_p => '0', value => x"015b"),
    (address => x"866691e", write_p => '0', value => x"015c"),
    (address => x"8666920", write_p => '0', value => x"015d"),
    (address => x"8666922", write_p => '0', value => x"015e"),
    (address => x"8666924", write_p => '0', value => x"015f"),
    (address => x"8666926", write_p => '0', value => x"0160"),
    (address => x"8666928", write_p => '0', value => x"0161"),
    (address => x"866692a", write_p => '0', value => x"0162"),
    (address => x"866692c", write_p => '0', value => x"0163"),
    (address => x"866692e", write_p => '0', value => x"0164"),
    (address => x"8666930", write_p => '0', value => x"0165"),
    (address => x"8666932", write_p => '0', value => x"0166"),
    (address => x"8666934", write_p => '0', value => x"0167"),
    (address => x"8666936", write_p => '0', value => x"0168"),
    (address => x"8666938", write_p => '0', value => x"0169"),
    (address => x"866693a", write_p => '0', value => x"016a"),
    (address => x"866693c", write_p => '0', value => x"016b"),
    (address => x"866693e", write_p => '0', value => x"016c"),
    (address => x"8666940", write_p => '0', value => x"016d"),
    (address => x"8666942", write_p => '0', value => x"016e"),
    (address => x"8666944", write_p => '0', value => x"016f"),
    (address => x"8666946", write_p => '0', value => x"0170"),
    (address => x"8666948", write_p => '0', value => x"0171"),
    (address => x"866694a", write_p => '0', value => x"0172"),
    (address => x"866694c", write_p => '0', value => x"0173"),
    (address => x"866694e", write_p => '0', value => x"0174"),
    (address => x"8666950", write_p => '0', value => x"0175"),
    (address => x"8666952", write_p => '0', value => x"0176"),
    (address => x"8666954", write_p => '0', value => x"0177"),
    (address => x"8666956", write_p => '0', value => x"0178"),
    (address => x"8666958", write_p => '0', value => x"0179"),
    (address => x"866695a", write_p => '0', value => x"017a"),
    (address => x"866695c", write_p => '0', value => x"017b"),
    (address => x"866695e", write_p => '0', value => x"017c"),
    (address => x"8666960", write_p => '0', value => x"017d"),
    (address => x"8666962", write_p => '0', value => x"017e"),
    (address => x"8666964", write_p => '0', value => x"017f"),
    (address => x"8666966", write_p => '0', value => x"0180"),
    (address => x"8666968", write_p => '0', value => x"0181"),
    (address => x"866696a", write_p => '0', value => x"0182"),
    (address => x"866696c", write_p => '0', value => x"0183"),
    (address => x"866696e", write_p => '0', value => x"0184"),
    (address => x"8666970", write_p => '0', value => x"0185"),
    (address => x"8666972", write_p => '0', value => x"0186"),
    (address => x"8666974", write_p => '0', value => x"0187"),
    (address => x"8666976", write_p => '0', value => x"0188"),
    (address => x"8666978", write_p => '0', value => x"0189"),
    (address => x"866697a", write_p => '0', value => x"018a"),
    (address => x"866697c", write_p => '0', value => x"018b"),
    (address => x"866697e", write_p => '0', value => x"018c"),
    (address => x"8666980", write_p => '0', value => x"018d"),
    (address => x"8666982", write_p => '0', value => x"018e"),
    (address => x"8666984", write_p => '0', value => x"018f"),
    (address => x"8666986", write_p => '0', value => x"0190"),
    (address => x"8666988", write_p => '0', value => x"0191"),
    (address => x"866698a", write_p => '0', value => x"0192"),
    (address => x"866698c", write_p => '0', value => x"0193"),
    (address => x"866698e", write_p => '0', value => x"0194"),
    (address => x"8666990", write_p => '0', value => x"0195"),
    (address => x"8666992", write_p => '0', value => x"0196"),
    (address => x"8666994", write_p => '0', value => x"0197"),
    (address => x"8666996", write_p => '0', value => x"0198"),
    (address => x"8666998", write_p => '0', value => x"0199"),
    (address => x"866699a", write_p => '0', value => x"019a"),
    (address => x"866699c", write_p => '0', value => x"019b"),
    (address => x"866699e", write_p => '0', value => x"019c"),
    (address => x"86669a0", write_p => '0', value => x"019d"),
    (address => x"86669a2", write_p => '0', value => x"019e"),
    (address => x"86669a4", write_p => '0', value => x"019f"),
    (address => x"86669a6", write_p => '0', value => x"01a0"),
    (address => x"86669a8", write_p => '0', value => x"01a1"),
    (address => x"86669aa", write_p => '0', value => x"01a2"),
    (address => x"86669ac", write_p => '0', value => x"01a3"),
    (address => x"86669ae", write_p => '0', value => x"01a4"),
    (address => x"86669b0", write_p => '0', value => x"01a5"),
    (address => x"86669b2", write_p => '0', value => x"01a6"),
    (address => x"86669b4", write_p => '0', value => x"01a7"),
    (address => x"86669b6", write_p => '0', value => x"01a8"),
    (address => x"86669b8", write_p => '0', value => x"01a9"),
    (address => x"86669ba", write_p => '0', value => x"01aa"),
    (address => x"86669bc", write_p => '0', value => x"01ab"),
    (address => x"86669be", write_p => '0', value => x"01ac"),
    (address => x"86669c0", write_p => '0', value => x"01ad"),
    (address => x"86669c2", write_p => '0', value => x"01ae"),
    (address => x"86669c4", write_p => '0', value => x"01af"),
    (address => x"86669c6", write_p => '0', value => x"01b0"),
    (address => x"86669c8", write_p => '0', value => x"01b1"),
    (address => x"86669ca", write_p => '0', value => x"01b2"),
    (address => x"86669cc", write_p => '0', value => x"01b3"),
    (address => x"86669ce", write_p => '0', value => x"01b4"),
    (address => x"86669d0", write_p => '0', value => x"01b5"),
    (address => x"86669d2", write_p => '0', value => x"01b6"),
    (address => x"86669d4", write_p => '0', value => x"01b7"),
    (address => x"86669d6", write_p => '0', value => x"01b8"),
    (address => x"86669d8", write_p => '0', value => x"01b9"),
    (address => x"86669da", write_p => '0', value => x"01ba"),
    (address => x"86669dc", write_p => '0', value => x"01bb"),
    (address => x"86669de", write_p => '0', value => x"01bc"),
    (address => x"86669e0", write_p => '0', value => x"01bd"),
    (address => x"86669e2", write_p => '0', value => x"01be"),
    (address => x"86669e4", write_p => '0', value => x"01bf"),
    (address => x"86669e6", write_p => '0', value => x"01c0"),
    (address => x"86669e8", write_p => '0', value => x"01c1"),
    (address => x"86669ea", write_p => '0', value => x"01c2"),
    (address => x"86669ec", write_p => '0', value => x"01c3"),
    (address => x"86669ee", write_p => '0', value => x"01c4"),
    (address => x"86669f0", write_p => '0', value => x"01c5"),
    (address => x"86669f2", write_p => '0', value => x"01c6"),
    (address => x"86669f4", write_p => '0', value => x"01c7"),
    (address => x"86669f6", write_p => '0', value => x"01c8"),
    (address => x"86669f8", write_p => '0', value => x"01c9"),
    (address => x"86669fa", write_p => '0', value => x"01ca"),
    (address => x"86669fc", write_p => '0', value => x"01cb"),
    (address => x"86669fe", write_p => '0', value => x"01cc"),
    (address => x"8666a00", write_p => '0', value => x"01cd"),
    (address => x"8666a02", write_p => '0', value => x"01ce"),
    (address => x"8666a04", write_p => '0', value => x"01cf"),
    (address => x"8666a06", write_p => '0', value => x"01d0"),
    (address => x"8666a08", write_p => '0', value => x"01d1"),
    (address => x"8666a0a", write_p => '0', value => x"01d2"),
    (address => x"8666a0c", write_p => '0', value => x"01d3"),
    (address => x"8666a0e", write_p => '0', value => x"01d4"),
    (address => x"8666a10", write_p => '0', value => x"01d5"),
    (address => x"8666a12", write_p => '0', value => x"01d6"),
    (address => x"8666a14", write_p => '0', value => x"01d7"),
    (address => x"8666a16", write_p => '0', value => x"01d8"),
    (address => x"8666a18", write_p => '0', value => x"01d9"),
    (address => x"8666a1a", write_p => '0', value => x"01da"),
    (address => x"8666a1c", write_p => '0', value => x"01db"),
    (address => x"8666a1e", write_p => '0', value => x"01dc"),
    (address => x"8666a20", write_p => '0', value => x"01dd"),
    (address => x"8666a22", write_p => '0', value => x"01de"),
    (address => x"8666a24", write_p => '0', value => x"01df"),
    (address => x"8666a26", write_p => '0', value => x"01e0"),
    (address => x"8666a28", write_p => '0', value => x"01e1"),
    (address => x"8666a2a", write_p => '0', value => x"01e2"),
    (address => x"8666a2c", write_p => '0', value => x"01e3"),
    (address => x"8666a2e", write_p => '0', value => x"01e4"),
    (address => x"8666a30", write_p => '0', value => x"01e5"),
    (address => x"8666a32", write_p => '0', value => x"01e6"),
    (address => x"8666a34", write_p => '0', value => x"01e7"),
    (address => x"8666a36", write_p => '0', value => x"01e8"),
    (address => x"8666a38", write_p => '0', value => x"01e9"),
    (address => x"8666a3a", write_p => '0', value => x"01ea"),
    (address => x"8666a3c", write_p => '0', value => x"01eb"),
    (address => x"8666a3e", write_p => '0', value => x"01ec"),
    (address => x"8666a40", write_p => '0', value => x"01ed"),
    (address => x"8666a42", write_p => '0', value => x"01ee"),
    (address => x"8666a44", write_p => '0', value => x"01ef"),
    (address => x"8666a46", write_p => '0', value => x"01f0"),
    (address => x"8666a48", write_p => '0', value => x"01f1"),
    (address => x"8666a4a", write_p => '0', value => x"01f2"),
    (address => x"8666a4c", write_p => '0', value => x"01f3"),
    (address => x"8666a4e", write_p => '0', value => x"01f4"),
    (address => x"8666a50", write_p => '0', value => x"01f5"),
    (address => x"8666a52", write_p => '0', value => x"01f6"),
    (address => x"8666a54", write_p => '0', value => x"01f7"),
    (address => x"8666a56", write_p => '0', value => x"01f8"),
    (address => x"8666a58", write_p => '0', value => x"01f9"),
    (address => x"8666a5a", write_p => '0', value => x"01fa"),
    (address => x"8666a5c", write_p => '0', value => x"01fb"),
    (address => x"8666a5e", write_p => '0', value => x"01fc"),
    (address => x"8666a60", write_p => '0', value => x"01fd"),
    (address => x"8666a62", write_p => '0', value => x"01fe"),
    (address => x"8666a64", write_p => '0', value => x"01ff"),
    (address => x"8666a66", write_p => '0', value => x"0200"),
    (address => x"8666a68", write_p => '0', value => x"0201"),
    (address => x"8666a6a", write_p => '0', value => x"0202"),
    (address => x"8666a6c", write_p => '0', value => x"0203"),
    (address => x"8666a6e", write_p => '0', value => x"0204"),
    (address => x"8666a70", write_p => '0', value => x"0205"),
    (address => x"8666a72", write_p => '0', value => x"0206"),
    (address => x"8666a74", write_p => '0', value => x"0207"),
    (address => x"8666a76", write_p => '0', value => x"0208"),
    (address => x"8666a78", write_p => '0', value => x"0209"),
    (address => x"8666a7a", write_p => '0', value => x"020a"),
    (address => x"8666a7c", write_p => '0', value => x"020b"),
    (address => x"8666a7e", write_p => '0', value => x"020c"),
    (address => x"8666a80", write_p => '0', value => x"020d"),
    (address => x"8666a82", write_p => '0', value => x"020e"),
    (address => x"8666a84", write_p => '0', value => x"020f"),
    (address => x"8666a86", write_p => '0', value => x"0210"),
    (address => x"8666a88", write_p => '0', value => x"0211"),
    (address => x"8666a8a", write_p => '0', value => x"0212"),
    (address => x"8666a8c", write_p => '0', value => x"0213"),
    (address => x"8666a8e", write_p => '0', value => x"0214"),
    (address => x"8666a90", write_p => '0', value => x"0215"),
    (address => x"8666a92", write_p => '0', value => x"0216"),
    (address => x"8666a94", write_p => '0', value => x"0217"),
    (address => x"8666a96", write_p => '0', value => x"0218"),
    (address => x"8666a98", write_p => '0', value => x"0219"),
    (address => x"8666a9a", write_p => '0', value => x"021a"),
    (address => x"8666a9c", write_p => '0', value => x"021b"),
    (address => x"8666a9e", write_p => '0', value => x"021c"),
    (address => x"8666aa0", write_p => '0', value => x"021d"),
    (address => x"8666aa2", write_p => '0', value => x"021e"),
    (address => x"8666aa4", write_p => '0', value => x"021f"),
    (address => x"8666aa6", write_p => '0', value => x"0220"),
    (address => x"8666aa8", write_p => '0', value => x"0221"),
    (address => x"8666aaa", write_p => '0', value => x"0222"),
    (address => x"8666aac", write_p => '0', value => x"0223"),
    (address => x"8666aae", write_p => '0', value => x"0224"),
    (address => x"8666ab0", write_p => '0', value => x"0225"),
    (address => x"8666ab2", write_p => '0', value => x"0226"),
    (address => x"8666ab4", write_p => '0', value => x"0227"),
    (address => x"8666ab6", write_p => '0', value => x"0228"),
    (address => x"8666ab8", write_p => '0', value => x"0229"),
    (address => x"8666aba", write_p => '0', value => x"022a"),
    (address => x"8666abc", write_p => '0', value => x"022b"),
    (address => x"8666abe", write_p => '0', value => x"022c"),
    (address => x"8666ac0", write_p => '0', value => x"022d"),
    (address => x"8666ac2", write_p => '0', value => x"022e"),
    (address => x"8666ac4", write_p => '0', value => x"022f"),
    (address => x"8666ac6", write_p => '0', value => x"0230"),
    (address => x"8666ac8", write_p => '0', value => x"0231"),
    (address => x"8666aca", write_p => '0', value => x"0232"),
    (address => x"8666acc", write_p => '0', value => x"0233"),
    (address => x"8666ace", write_p => '0', value => x"0234"),
    (address => x"8666ad0", write_p => '0', value => x"0235"),
    (address => x"8666ad2", write_p => '0', value => x"0236"),
    (address => x"8666ad4", write_p => '0', value => x"0237"),
    (address => x"8666ad6", write_p => '0', value => x"0238"),
    (address => x"8666ad8", write_p => '0', value => x"0239"),
    (address => x"8666ada", write_p => '0', value => x"023a"),
    (address => x"8666adc", write_p => '0', value => x"023b"),
    (address => x"8666ade", write_p => '0', value => x"023c"),
    (address => x"8666ae0", write_p => '0', value => x"023d"),
    (address => x"8666ae2", write_p => '0', value => x"023e"),
    (address => x"8666ae4", write_p => '0', value => x"023f"),
    (address => x"8666ae6", write_p => '0', value => x"0240"),
    (address => x"8666ae8", write_p => '0', value => x"0241"),
    (address => x"8666aea", write_p => '0', value => x"0242"),
    (address => x"8666aec", write_p => '0', value => x"0243"),
    (address => x"8666aee", write_p => '0', value => x"0244"),
    (address => x"8666af0", write_p => '0', value => x"0245"),
    (address => x"8666af2", write_p => '0', value => x"0246"),
    (address => x"8666af4", write_p => '0', value => x"0247"),
    (address => x"8666af6", write_p => '0', value => x"0248"),
    (address => x"8666af8", write_p => '0', value => x"0249"),
    (address => x"8666afa", write_p => '0', value => x"024a"),
    (address => x"8666afc", write_p => '0', value => x"024b"),
    (address => x"8666afe", write_p => '0', value => x"024c"),
    (address => x"8666b00", write_p => '0', value => x"024d"),
    (address => x"8666b02", write_p => '0', value => x"024e"),
    (address => x"8666b04", write_p => '0', value => x"024f"),
    (address => x"8666b06", write_p => '0', value => x"0250"),
    (address => x"8666b08", write_p => '0', value => x"0251"),
    (address => x"8666b0a", write_p => '0', value => x"0252"),
    (address => x"8666b0c", write_p => '0', value => x"0253"),
    (address => x"8666b0e", write_p => '0', value => x"0254"),
    (address => x"8666b10", write_p => '0', value => x"0255"),
    (address => x"8666b12", write_p => '0', value => x"0256"),
    (address => x"8666b14", write_p => '0', value => x"0257"),
    (address => x"8666b16", write_p => '0', value => x"0258"),
    (address => x"8666b18", write_p => '0', value => x"0259"),
    (address => x"8666b1a", write_p => '0', value => x"025a"),
    (address => x"8666b1c", write_p => '0', value => x"025b"),
    (address => x"8666b1e", write_p => '0', value => x"025c"),
    (address => x"8666b20", write_p => '0', value => x"025d"),
    (address => x"8666b22", write_p => '0', value => x"025e"),
    (address => x"8666b24", write_p => '0', value => x"025f"),
    (address => x"8666b26", write_p => '0', value => x"0260"),
    (address => x"8666b28", write_p => '0', value => x"0261"),
    (address => x"8666b2a", write_p => '0', value => x"0262"),
    (address => x"8666b2c", write_p => '0', value => x"0263"),
    (address => x"8666b2e", write_p => '0', value => x"0264"),
    (address => x"8666b30", write_p => '0', value => x"0265"),
    (address => x"8666b32", write_p => '0', value => x"0266"),
    (address => x"8666b34", write_p => '0', value => x"0267"),
    (address => x"8666b36", write_p => '0', value => x"0268"),
    (address => x"8666b38", write_p => '0', value => x"0269"),
    (address => x"8666b3a", write_p => '0', value => x"026a"),
    (address => x"8666b3c", write_p => '0', value => x"026b"),
    (address => x"8666b3e", write_p => '0', value => x"026c"),
    (address => x"8666b40", write_p => '0', value => x"026d"),
    (address => x"8666b42", write_p => '0', value => x"026e"),
    (address => x"8666b44", write_p => '0', value => x"026f"),
    (address => x"8666b46", write_p => '0', value => x"0270"),
    (address => x"8666b48", write_p => '0', value => x"0271"),
    (address => x"8666b4a", write_p => '0', value => x"0272"),
    (address => x"8666b4c", write_p => '0', value => x"0273"),
    (address => x"8666b4e", write_p => '0', value => x"0274"),
    (address => x"8666b50", write_p => '0', value => x"0275"),
    (address => x"8666b52", write_p => '0', value => x"0276"),
    (address => x"8666b54", write_p => '0', value => x"0277"),
    (address => x"8666b56", write_p => '0', value => x"0278"),
    (address => x"8666b58", write_p => '0', value => x"0279"),
    (address => x"8666b5a", write_p => '0', value => x"027a"),
    (address => x"8666b5c", write_p => '0', value => x"027b"),
    (address => x"8666b5e", write_p => '0', value => x"027c"),
    (address => x"8666b60", write_p => '0', value => x"027d"),
    (address => x"8666b62", write_p => '0', value => x"027e"),
    (address => x"8666b64", write_p => '0', value => x"027f"),
    (address => x"8666b66", write_p => '0', value => x"0280"),
    (address => x"8666b68", write_p => '0', value => x"0281"),
    (address => x"8666b6a", write_p => '0', value => x"0282"),
    (address => x"8666b6c", write_p => '0', value => x"0283"),
    (address => x"8666b6e", write_p => '0', value => x"0284"),
    (address => x"8666b70", write_p => '0', value => x"0285"),
    (address => x"8666b72", write_p => '0', value => x"0286"),
    (address => x"8666b74", write_p => '0', value => x"0287"),
    (address => x"8666b76", write_p => '0', value => x"0288"),
    (address => x"8666b78", write_p => '0', value => x"0289"),
    (address => x"8666b7a", write_p => '0', value => x"028a"),
    (address => x"8666b7c", write_p => '0', value => x"028b"),
    (address => x"8666b7e", write_p => '0', value => x"028c"),
    (address => x"8666b80", write_p => '0', value => x"028d"),
    (address => x"8666b82", write_p => '0', value => x"028e"),
    (address => x"8666b84", write_p => '0', value => x"028f"),
    (address => x"8666b86", write_p => '0', value => x"0290"),
    (address => x"8666b88", write_p => '0', value => x"0291"),
    (address => x"8666b8a", write_p => '0', value => x"0292"),
    (address => x"8666b8c", write_p => '0', value => x"0293"),
    (address => x"8666b8e", write_p => '0', value => x"0294"),
    (address => x"8666b90", write_p => '0', value => x"0295"),
    (address => x"8666b92", write_p => '0', value => x"0296"),
    (address => x"8666b94", write_p => '0', value => x"0297"),
    (address => x"8666b96", write_p => '0', value => x"0298"),
    (address => x"8666b98", write_p => '0', value => x"0299"),
    (address => x"8666b9a", write_p => '0', value => x"029a"),
    (address => x"8666b9c", write_p => '0', value => x"029b"),
    (address => x"8666b9e", write_p => '0', value => x"029c"),
    (address => x"8666ba0", write_p => '0', value => x"029d"),
    (address => x"8666ba2", write_p => '0', value => x"029e"),
    (address => x"8666ba4", write_p => '0', value => x"029f"),
    (address => x"8666ba6", write_p => '0', value => x"02a0"),
    (address => x"8666ba8", write_p => '0', value => x"02a1"),
    (address => x"8666baa", write_p => '0', value => x"02a2"),
    (address => x"8666bac", write_p => '0', value => x"02a3"),
    (address => x"8666bae", write_p => '0', value => x"02a4"),
    (address => x"8666bb0", write_p => '0', value => x"02a5"),
    (address => x"8666bb2", write_p => '0', value => x"02a6"),
    (address => x"8666bb4", write_p => '0', value => x"02a7"),
    (address => x"8666bb6", write_p => '0', value => x"02a8"),
    (address => x"8666bb8", write_p => '0', value => x"02a9"),
    (address => x"8666bba", write_p => '0', value => x"02aa"),
    (address => x"8666bbc", write_p => '0', value => x"02ab"),
    (address => x"8666bbe", write_p => '0', value => x"02ac"),
    (address => x"8666bc0", write_p => '0', value => x"02ad"),
    (address => x"8666bc2", write_p => '0', value => x"02ae"),
    (address => x"8666bc4", write_p => '0', value => x"02af"),
    (address => x"8666bc6", write_p => '0', value => x"02b0"),
    (address => x"8666bc8", write_p => '0', value => x"02b1"),
    (address => x"8666bca", write_p => '0', value => x"02b2"),
    (address => x"8666bcc", write_p => '0', value => x"02b3"),
    (address => x"8666bce", write_p => '0', value => x"02b4"),
    (address => x"8666bd0", write_p => '0', value => x"02b5"),
    (address => x"8666bd2", write_p => '0', value => x"02b6"),
    (address => x"8666bd4", write_p => '0', value => x"02b7"),
    (address => x"8666bd6", write_p => '0', value => x"02b8"),
    (address => x"8666bd8", write_p => '0', value => x"02b9"),
    (address => x"8666bda", write_p => '0', value => x"02ba"),
    (address => x"8666bdc", write_p => '0', value => x"02bb"),
    (address => x"8666bde", write_p => '0', value => x"02bc"),
    (address => x"8666be0", write_p => '0', value => x"02bd"),
    (address => x"8666be2", write_p => '0', value => x"02be"),
    (address => x"8666be4", write_p => '0', value => x"02bf"),
    (address => x"8666be6", write_p => '0', value => x"02c0"),
    (address => x"8666be8", write_p => '0', value => x"02c1"),
    (address => x"8666bea", write_p => '0', value => x"02c2"),
    (address => x"8666bec", write_p => '0', value => x"02c3"),
    (address => x"8666bee", write_p => '0', value => x"02c4"),
    (address => x"8666bf0", write_p => '0', value => x"02c5"),
    (address => x"8666bf2", write_p => '0', value => x"02c6"),
    (address => x"8666bf4", write_p => '0', value => x"02c7"),
    (address => x"8666bf6", write_p => '0', value => x"02c8"),
    (address => x"8666bf8", write_p => '0', value => x"02c9"),
    (address => x"8666bfa", write_p => '0', value => x"02ca"),
    (address => x"8666bfc", write_p => '0', value => x"02cb"),
    (address => x"8666bfe", write_p => '0', value => x"02cc"),
    (address => x"8666c00", write_p => '0', value => x"02cd"),
    (address => x"8666c02", write_p => '0', value => x"02ce"),
    (address => x"8666c04", write_p => '0', value => x"02cf"),
    (address => x"8666c06", write_p => '0', value => x"02d0"),
    (address => x"8666c08", write_p => '0', value => x"02d1"),
    (address => x"8666c0a", write_p => '0', value => x"02d2"),
    (address => x"8666c0c", write_p => '0', value => x"02d3"),
    (address => x"8666c0e", write_p => '0', value => x"02d4"),
    (address => x"8666c10", write_p => '0', value => x"02d5"),
    (address => x"8666c12", write_p => '0', value => x"02d6"),
    (address => x"8666c14", write_p => '0', value => x"02d7"),
    (address => x"8666c16", write_p => '0', value => x"02d8"),
    (address => x"8666c18", write_p => '0', value => x"02d9"),
    (address => x"8666c1a", write_p => '0', value => x"02da"),
    (address => x"8666c1c", write_p => '0', value => x"02db"),
    (address => x"8666c1e", write_p => '0', value => x"02dc"),
    (address => x"8666c20", write_p => '0', value => x"02dd"),
    (address => x"8666c22", write_p => '0', value => x"02de"),
    (address => x"8666c24", write_p => '0', value => x"02df"),
    (address => x"8666c26", write_p => '0', value => x"02e0"),
    (address => x"8666c28", write_p => '0', value => x"02e1"),
    (address => x"8666c2a", write_p => '0', value => x"02e2"),
    (address => x"8666c2c", write_p => '0', value => x"02e3"),
    (address => x"8666c2e", write_p => '0', value => x"02e4"),
    (address => x"8666c30", write_p => '0', value => x"02e5"),
    (address => x"8666c32", write_p => '0', value => x"02e6"),
    (address => x"8666c34", write_p => '0', value => x"02e7"),
    (address => x"8666c36", write_p => '0', value => x"02e8"),
    (address => x"8666c38", write_p => '0', value => x"02e9"),
    (address => x"8666c3a", write_p => '0', value => x"02ea"),
    (address => x"8666c3c", write_p => '0', value => x"02eb"),
    (address => x"8666c3e", write_p => '0', value => x"02ec"),
    (address => x"8666c40", write_p => '0', value => x"02ed"),
    (address => x"8666c42", write_p => '0', value => x"02ee"),
    (address => x"8666c44", write_p => '0', value => x"02ef"),
    (address => x"8666c46", write_p => '0', value => x"02f0"),
    (address => x"8666c48", write_p => '0', value => x"02f1"),
    (address => x"8666c4a", write_p => '0', value => x"02f2"),
    (address => x"8666c4c", write_p => '0', value => x"02f3"),
    (address => x"8666c4e", write_p => '0', value => x"02f4"),
    (address => x"8666c50", write_p => '0', value => x"02f5"),
    (address => x"8666c52", write_p => '0', value => x"02f6"),
    (address => x"8666c54", write_p => '0', value => x"02f7"),
    (address => x"8666c56", write_p => '0', value => x"02f8"),
    (address => x"8666c58", write_p => '0', value => x"02f9"),
    (address => x"8666c5a", write_p => '0', value => x"02fa"),
    (address => x"8666c5c", write_p => '0', value => x"02fb"),
    (address => x"8666c5e", write_p => '0', value => x"02fc"),
    (address => x"8666c60", write_p => '0', value => x"02fd"),
    (address => x"8666c62", write_p => '0', value => x"02fe"),
    (address => x"8666c64", write_p => '0', value => x"02ff"),
    
    
    
    others => ( address => x"FFFFFFF", write_p => '0', value => x"0000")
    );

  -- Wait initially to allow hyperram to reset and set config register
  signal idle_wait : std_logic := '0';
  
  signal expect_value : std_logic := '0';
  signal expected_value : unsigned(15 downto 0) := x"0000";

  signal viciv_addr : unsigned(18 downto 3) := (others => '0');
  signal viciv_request_toggle : std_logic := '0';
  signal viciv_data : unsigned(7 downto 0) := x"00";
  signal viciv_data_strobe : std_logic := '0';
  signal pixel_counter : unsigned(31 downto 0) := to_unsigned(0,32);
  
begin

--  reconfig1: entity work.reconfig
--    port map ( clock => clock163,
--               trigger_reconfigure => '0',
--               reconfigure_address => (others => '0'));
  
  hyperram0: entity work.hyperram
    generic map ( in_simulation => true )
    port map (
      pixelclock => pixelclock,
      clock163 => clock163,
      clock325 => clock325,
      address => expansionram_address,
      wdata => expansionram_wdata(7 downto 0),
      wdata_hi => expansionram_wdata(15 downto 8),
      wen_hi => '1',
      wen_lo => '1',
      read_request => expansionram_read,
      write_request => expansionram_write,
      rdata_16en => '1',
      rdata => expansionram_rdata(7 downto 0),
      rdata_hi =>  expansionram_rdata(15 downto 8),
      data_ready_strobe => expansionram_data_ready_strobe,
      busy => expansionram_busy,

      current_cache_line => current_cache_line,
      current_cache_line_address => current_cache_line_address,
      current_cache_line_valid => current_cache_line_valid,
      expansionram_current_cache_line_next_toggle  => expansionram_current_cache_line_next_toggle,

      viciv_addr => viciv_addr,
      viciv_request_toggle => viciv_request_toggle,
      viciv_data_out => viciv_data,
      viciv_data_strobe => viciv_data_strobe,
      
      hr_d => hr_d,
      hr_rwds => hr_rwds,
      hr_reset => hr_reset,
      hr_clk_n => hr_clk_n,
      hr_clk_p => hr_clk_p,
      hr_cs0 => hr_cs0,

      hr2_d => hr2_d,
      hr2_rwds => hr2_rwds,
      hr2_reset => hr2_reset,
      hr2_clk_n => hr2_clk_n,
      hr2_clk_p => hr2_clk_p,
      hr_cs1 => hr2_cs0
      
      );

  fakehyper0: entity work.s27kl0641
    generic map (
      id => "$8000000",
      tdevice_vcs => 5 ns,
      timingmodel => "S27KL0641DABHI000"
      )
    port map (
      DQ7 => hr_d(7),
      DQ6 => hr_d(6),
      DQ5 => hr_d(5),
      DQ4 => hr_d(4),
      DQ3 => hr_d(3),
      DQ2 => hr_d(2),
      DQ1 => hr_d(1),
      DQ0 => hr_d(0),

      CSNeg => hr_cs0,
      CK => hr_clk_p,
      RESETneg => hr_reset,
      RWDS => hr_rwds
      );
  

  fakehyper1: entity work.s27kl0641
    generic map (
      id => "$8800000",
      tdevice_vcs => 5 ns,
      timingmodel => "S27KL0641DABHI000"
      )
    port map (
      DQ7 => hr2_d(7),
      DQ6 => hr2_d(6),
      DQ5 => hr2_d(5),
      DQ4 => hr2_d(4),
      DQ3 => hr2_d(3),
      DQ2 => hr2_d(2),
      DQ1 => hr2_d(1),
      DQ0 => hr2_d(0),

      CSNeg => hr2_cs0,
      CK => hr2_clk_p,
      RESETneg => hr2_reset,
      RWDS => hr2_rwds
      );
  
  process(hr_cs0, hr_clk_p, hr_reset, hr_rwds, hr_d,
          hr2_cs0, hr2_clk_p, hr2_reset, hr2_rwds, hr2_d
          ) is
  begin
    if true then
      report
        "hr_cs0 = " & std_logic'image(hr_cs0) & ", " &
        "hr_clk_p = " & std_logic'image(hr_clk_p) & ", " &
        "hr_reset = " & std_logic'image(hr_reset) & ", " &
        "hr_rwds = " & std_logic'image(hr_rwds) & ", " &
        "hr_d = " & std_logic'image(hr_d(0))
        & std_logic'image(hr_d(1))
        & std_logic'image(hr_d(2))
        & std_logic'image(hr_d(3))
        & std_logic'image(hr_d(4))
        & std_logic'image(hr_d(5))
        & std_logic'image(hr_d(6))
        & std_logic'image(hr_d(7))
        & ".";
      report
        "hr2_cs0 = " & std_logic'image(hr2_cs0) & ", " &
        "hr2_clk_p = " & std_logic'image(hr2_clk_p) & ", " &
        "hr2_reset = " & std_logic'image(hr2_reset) & ", " &
        "hr2_rwds = " & std_logic'image(hr2_rwds) & ", " &
        "hr2_d = " & std_logic'image(hr2_d(0))
        & std_logic'image(hr2_d(1))
        & std_logic'image(hr2_d(2))
        & std_logic'image(hr2_d(3))
        & std_logic'image(hr2_d(4))
        & std_logic'image(hr2_d(5))
        & std_logic'image(hr2_d(6))
        & std_logic'image(hr2_d(7))
        & ".";
    end if;
  end process;

  process (pixelclock) is
  begin
    if false and rising_edge(pixelclock) then
      pixel_counter <= pixel_counter + 1;
      if (pixel_counter(9 downto 0) = to_unsigned(0,10)) then
        report "VIC: Dispatching pixel data request";
        viciv_request_toggle <= pixel_counter(10);
        viciv_addr <= pixel_counter(23 downto 8);
      end if;
      if viciv_data_strobe='1' then
        report "VIC: Received byte $" & to_hstring(viciv_data);
      end if;
    end if;
  end process;
  
  
  process (clock325) is
  begin
    if rising_edge(clock325) then
      current_time <= current_time + 3;
    end if;
  end process;
  
  process (pixelclock) is
  begin

    if rising_edge(pixelclock) then

      if true then
        report "expansionram_data_ready_strobe=" & std_logic'image(expansionram_data_ready_strobe) 
          & ", expansionram_busy=" & std_logic'image(expansionram_busy)
          & ", expansionram_read=" & std_logic'image(expansionram_read)
          & ", idle_wait=" & std_logic'image(idle_wait)
          & ", expect_value=" & std_logic'image(expect_value);
      end if;
      
      if expansionram_data_ready_strobe='1' then
        if expect_value = '1' then
          if expected_value = expansionram_rdata then
            report "DISPATCHER: Read correct value $" & to_hstring(expansionram_rdata)
              & " after " & integer'image(current_time - dispatch_time) & "ns.";
          else
            report "DISPATCHER: ERROR: Expected $" & to_hstring(expected_value) & ", but saw $" & to_hstring(expansionram_rdata)
              & " after " & integer'image(current_time - dispatch_time) & "ns.";            
          end if;
          dispatch_time <= current_time;
        end if;        
        expect_value <= '0';
        idle_wait <= '0';
      end if;

      expansionram_write <= '0';
      expansionram_read <= '0';

      if expansionram_busy='1' then
        idle_wait <= '0';
      else
        if expect_value = '0' and expansionram_busy='0' then

          if expansionram_busy = '0' and idle_wait='0' then

            if mem_jobs(cycles).address = x"FFFFFFF" then
              report "DISPATCHER: Total sequence was " & integer'image(current_time - start_time) & "ns "
                & "(mean " & integer'image(1+(current_time-start_time)/cycles) & "ns ).";
              cycles <= 0;
              start_time <= current_time;          
            else
              cycles <= cycles + 1;        
            end if;

            dispatch_time <= current_time;
            
            expansionram_address <= mem_jobs(cycles).address(26 downto 0);
            expansionram_write <= mem_jobs(cycles).write_p;
            expansionram_read <= not mem_jobs(cycles).write_p;
            expansionram_wdata <= mem_jobs(cycles).value;
            -- Only wait for memory reads?
            idle_wait <= not mem_jobs(cycles).write_p;

            if (mem_jobs(cycles).write_p='0') then
              -- Let reads finish serially
              -- (In the worst case, this can take quite a while)
              report "DISPATCHER: Reading from $" & to_hstring(mem_jobs(cycles).address) & ", expecting to see $"
                & to_hstring(mem_jobs(cycles).value);
              expect_value <= '1';
              expected_value <= mem_jobs(cycles).value;
            else
              report "DISPATCHER: Writing to $" & to_hstring(mem_jobs(cycles).address) & " <- $"
                & to_hstring(mem_jobs(cycles).value);
              expect_value <= '0';
              dispatch_time <= current_time;
            end if;

            if start_time = 0 then
              start_time <= current_time;
            end if;
          end if;
        end if;
      end if;
    end if;
    
  end process;

  process is
  begin
    
    clock325 <= '0';
    pixelclock <= '0';
    cpuclock <= '0';
    clock163 <= '0';

    report "tick";
    
    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;
    
    clock163 <= '1';

    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    pixelclock <= '1';
    clock163 <= '0';

    report "tick";   
    
    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    clock163 <= '1';

    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    pixelclock <= '0';
    cpuclock <= '1';
    clock163 <= '0';

    report "tick";    

    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    clock163 <= '1';

    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    pixelclock <= '1';
    clock163 <= '0';

    report "tick";
    
    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

    clock163 <= '1';

    clock325 <= '1';
    wait for 1.5 ns;
    clock325 <= '0';
    wait for 1.5 ns;

--    report "40MHz CPU clock cycle finished";
    
  end process;


end foo;
