
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity BLE_4 is
	port ( clk          : in  std_ulogic;
	       rst          : in  std_ulogic;
	       --------------------------------------------------
	       clk_app      : in  std_ulogic;
	       --------------------------------------------------
	       snap_in      : in  std_ulogic;
	       snap_out     : out std_ulogic;
	       snap_restore : in  std_ulogic;
	       --------------------------------------------------
	       config       : in  std_ulogic_vector(16 downto 0);
	       inputs       : in  std_ulogic_vector(3 downto 0);
	       output       : out std_ulogic);
end BLE_4;


architecture RTL of BLE_4 is

	signal reg_config : std_ulogic := '0';
	signal lut_config : std_ulogic_vector(15 downto 0) := (others => '0');
	signal lut_output : std_ulogic := '0';
	signal reg_output : std_ulogic := '0';

begin

	reg_config <= config(16);
	lut_config <= config(15 downto 0);

	lut_output <= lut_config(to_integer(unsigned(inputs)));

	process(clk)
	begin
		if rising_edge(clk) then
			if rst = '1' then
				reg_output <= '0';
			elsif snap_restore = '1' then
				reg_output <= snap_in;
			elsif clk_app = '1' then
				reg_output <= lut_output;
			end if;
		end if;
	end process;

	snap_out <= reg_output;

	output <= reg_output when reg_config = '1' else lut_output;

end RTL;


--------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity CLB_clb_N4K4I10O4 is
	port ( clk          : in  std_ulogic;
	       rst          : in  std_ulogic;
	       --------------------------------------------------
	       clk_app      : in  std_ulogic;
	       --------------------------------------------------
	       snap_in      : in  std_ulogic_vector(3 downto 0);
	       snap_out     : out std_ulogic_vector(3 downto 0);
	       snap_restore : in  std_ulogic;
	       --------------------------------------------------
	       config       : in  std_ulogic_vector(131 downto 0);
	       inputs       : in  std_ulogic_vector(9 downto 0);
	       outputs      : out std_ulogic_vector(3 downto 0));
end CLB_clb_N4K4I10O4;


architecture RTL of CLB_clb_N4K4I10O4 is

	signal outputs_int          : std_ulogic_vector(3 downto 0) := (others => '0');

	signal crossbar_inputs      : std_ulogic_vector(15 downto 0) := (others => '0');
	signal crossbar_outputs     : std_ulogic_vector(15 downto 0) := (others => '0');

	signal crossbar_selector_00 : integer range 0 to 15 := 0;
	signal crossbar_selector_01 : integer range 0 to 15 := 0;
	signal crossbar_selector_02 : integer range 0 to 15 := 0;
	signal crossbar_selector_03 : integer range 0 to 15 := 0;
	signal crossbar_selector_04 : integer range 0 to 15 := 0;
	signal crossbar_selector_05 : integer range 0 to 15 := 0;
	signal crossbar_selector_06 : integer range 0 to 15 := 0;
	signal crossbar_selector_07 : integer range 0 to 15 := 0;
	signal crossbar_selector_08 : integer range 0 to 15 := 0;
	signal crossbar_selector_09 : integer range 0 to 15 := 0;
	signal crossbar_selector_10 : integer range 0 to 15 := 0;
	signal crossbar_selector_11 : integer range 0 to 15 := 0;
	signal crossbar_selector_12 : integer range 0 to 15 := 0;
	signal crossbar_selector_13 : integer range 0 to 15 := 0;
	signal crossbar_selector_14 : integer range 0 to 15 := 0;
	signal crossbar_selector_15 : integer range 0 to 15 := 0;

begin

	crossbar_inputs <= "00" & outputs_int & inputs;

	crossbar_selector_00 <= to_integer(unsigned(config(71 downto 68)));
	crossbar_selector_01 <= to_integer(unsigned(config(75 downto 72)));
	crossbar_selector_02 <= to_integer(unsigned(config(79 downto 76)));
	crossbar_selector_03 <= to_integer(unsigned(config(83 downto 80)));
	crossbar_selector_04 <= to_integer(unsigned(config(87 downto 84)));
	crossbar_selector_05 <= to_integer(unsigned(config(91 downto 88)));
	crossbar_selector_06 <= to_integer(unsigned(config(95 downto 92)));
	crossbar_selector_07 <= to_integer(unsigned(config(99 downto 96)));
	crossbar_selector_08 <= to_integer(unsigned(config(103 downto 100)));
	crossbar_selector_09 <= to_integer(unsigned(config(107 downto 104)));
	crossbar_selector_10 <= to_integer(unsigned(config(111 downto 108)));
	crossbar_selector_11 <= to_integer(unsigned(config(115 downto 112)));
	crossbar_selector_12 <= to_integer(unsigned(config(119 downto 116)));
	crossbar_selector_13 <= to_integer(unsigned(config(123 downto 120)));
	crossbar_selector_14 <= to_integer(unsigned(config(127 downto 124)));
	crossbar_selector_15 <= to_integer(unsigned(config(131 downto 128)));

	-- Virtual Time Propagation Registers are placed between the CLB crossbar and BLE inputs --
	process(clk)
	begin
		if rising_edge(clk) then
			crossbar_outputs(0) <= crossbar_inputs(crossbar_selector_00);
			crossbar_outputs(1) <= crossbar_inputs(crossbar_selector_01);
			crossbar_outputs(2) <= crossbar_inputs(crossbar_selector_02);
			crossbar_outputs(3) <= crossbar_inputs(crossbar_selector_03);
			crossbar_outputs(4) <= crossbar_inputs(crossbar_selector_04);
			crossbar_outputs(5) <= crossbar_inputs(crossbar_selector_05);
			crossbar_outputs(6) <= crossbar_inputs(crossbar_selector_06);
			crossbar_outputs(7) <= crossbar_inputs(crossbar_selector_07);
			crossbar_outputs(8) <= crossbar_inputs(crossbar_selector_08);
			crossbar_outputs(9) <= crossbar_inputs(crossbar_selector_09);
			crossbar_outputs(10) <= crossbar_inputs(crossbar_selector_10);
			crossbar_outputs(11) <= crossbar_inputs(crossbar_selector_11);
			crossbar_outputs(12) <= crossbar_inputs(crossbar_selector_12);
			crossbar_outputs(13) <= crossbar_inputs(crossbar_selector_13);
			crossbar_outputs(14) <= crossbar_inputs(crossbar_selector_14);
			crossbar_outputs(15) <= crossbar_inputs(crossbar_selector_15);
		end if;
	end process;

	BLE4_0: entity work.BLE_4
	port map ( clk           => clk,
	           rst           => rst,
	           clk_app       => clk_app,
	           snap_in       => snap_in(0),
	           snap_out      => snap_out(0),
	           snap_restore  => snap_restore,
	           config        => config(16 downto 0),
	           inputs        => crossbar_outputs(3 downto 0),
	           output        => outputs_int(0));

	BLE4_1: entity work.BLE_4
	port map ( clk           => clk,
	           rst           => rst,
	           clk_app       => clk_app,
	           snap_in       => snap_in(1),
	           snap_out      => snap_out(1),
	           snap_restore  => snap_restore,
	           config        => config(33 downto 17),
	           inputs        => crossbar_outputs(7 downto 4),
	           output        => outputs_int(1));

	BLE4_2: entity work.BLE_4
	port map ( clk           => clk,
	           rst           => rst,
	           clk_app       => clk_app,
	           snap_in       => snap_in(2),
	           snap_out      => snap_out(2),
	           snap_restore  => snap_restore,
	           config        => config(50 downto 34),
	           inputs        => crossbar_outputs(11 downto 8),
	           output        => outputs_int(2));

	BLE4_3: entity work.BLE_4
	port map ( clk           => clk,
	           rst           => rst,
	           clk_app       => clk_app,
	           snap_in       => snap_in(3),
	           snap_out      => snap_out(3),
	           snap_restore  => snap_restore,
	           config        => config(67 downto 51),
	           inputs        => crossbar_outputs(15 downto 12),
	           output        => outputs_int(3));

	outputs <= outputs_int;

end RTL;


--------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_matrix is
	port ( clk          : in  std_ulogic;
	       rst          : in  std_ulogic;
	       --------------------------------------------------
	       clk_app      : in  std_ulogic;
	       --------------------------------------------------
	       config       : in  std_ulogic_vector(10951 downto 0);
	       --------------------------------------------------
	       snap_in      : in  std_ulogic_vector(191 downto 0);
	       snap_out     : out std_ulogic_vector(191 downto 0);
	       snap_restore : in  std_ulogic;
	       --------------------------------------------------
	       inputs       : in  std_ulogic_vector(55 downto 0);
	       outputs      : out std_ulogic_vector(55 downto 0));
end ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_matrix;


architecture RTL of ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_matrix is

	-- Output pins (for CLBs and IOs) --
	signal CLB_1_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_1_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_1_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_1_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_1_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_1_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_1_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_1_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_1_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_2_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_2_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_2_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_2_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_3_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_3_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_3_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_3_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_4_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_4_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_4_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_4_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_5_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_5_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_5_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_5_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_6_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_6_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_6_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_6_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_7_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_7_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_7_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_7_6_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_1_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_1_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_1_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_1_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_2_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_2_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_2_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_2_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_3_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_3_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_3_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_3_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_4_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_4_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_4_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_4_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_5_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_5_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_5_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_5_OUT_pin_3 : std_ulogic := '0';
	signal CLB_8_6_OUT_pin_0 : std_ulogic := '0';
	signal CLB_8_6_OUT_pin_1 : std_ulogic := '0';
	signal CLB_8_6_OUT_pin_2 : std_ulogic := '0';
	signal CLB_8_6_OUT_pin_3 : std_ulogic := '0';
	signal IO_0_1_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_1_OUT_pin_1  : std_ulogic := '0';
	signal IO_0_2_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_2_OUT_pin_1  : std_ulogic := '0';
	signal IO_0_3_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_3_OUT_pin_1  : std_ulogic := '0';
	signal IO_0_4_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_4_OUT_pin_1  : std_ulogic := '0';
	signal IO_0_5_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_5_OUT_pin_1  : std_ulogic := '0';
	signal IO_0_6_OUT_pin_0  : std_ulogic := '0';
	signal IO_0_6_OUT_pin_1  : std_ulogic := '0';
	signal IO_1_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_1_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_1_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_1_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_2_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_2_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_2_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_2_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_3_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_3_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_3_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_3_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_4_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_4_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_4_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_4_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_5_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_5_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_5_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_5_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_6_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_6_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_6_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_6_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_7_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_7_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_7_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_7_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_8_0_OUT_pin_0  : std_ulogic := '0';
	signal IO_8_0_OUT_pin_1  : std_ulogic := '0';
	signal IO_8_7_OUT_pin_0  : std_ulogic := '0';
	signal IO_8_7_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_1_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_1_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_2_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_2_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_3_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_3_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_4_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_4_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_5_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_5_OUT_pin_1  : std_ulogic := '0';
	signal IO_9_6_OUT_pin_0  : std_ulogic := '0';
	signal IO_9_6_OUT_pin_1  : std_ulogic := '0';

	-- Input pins (for CLBs and IOs) --
	signal CLB_1_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_1_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_2_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_3_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_4_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_5_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_6_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_7_6_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_1_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_2_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_3_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_4_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_5_IN_pin_9 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_0 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_1 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_2 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_3 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_4 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_5 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_6 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_7 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_8 : std_ulogic := '0';
	signal CLB_8_6_IN_pin_9 : std_ulogic := '0';
	signal IO_0_1_IN_pin_0  : std_ulogic := '0';
	signal IO_0_1_IN_pin_1  : std_ulogic := '0';
	signal IO_0_2_IN_pin_0  : std_ulogic := '0';
	signal IO_0_2_IN_pin_1  : std_ulogic := '0';
	signal IO_0_3_IN_pin_0  : std_ulogic := '0';
	signal IO_0_3_IN_pin_1  : std_ulogic := '0';
	signal IO_0_4_IN_pin_0  : std_ulogic := '0';
	signal IO_0_4_IN_pin_1  : std_ulogic := '0';
	signal IO_0_5_IN_pin_0  : std_ulogic := '0';
	signal IO_0_5_IN_pin_1  : std_ulogic := '0';
	signal IO_0_6_IN_pin_0  : std_ulogic := '0';
	signal IO_0_6_IN_pin_1  : std_ulogic := '0';
	signal IO_1_0_IN_pin_0  : std_ulogic := '0';
	signal IO_1_0_IN_pin_1  : std_ulogic := '0';
	signal IO_1_7_IN_pin_0  : std_ulogic := '0';
	signal IO_1_7_IN_pin_1  : std_ulogic := '0';
	signal IO_2_0_IN_pin_0  : std_ulogic := '0';
	signal IO_2_0_IN_pin_1  : std_ulogic := '0';
	signal IO_2_7_IN_pin_0  : std_ulogic := '0';
	signal IO_2_7_IN_pin_1  : std_ulogic := '0';
	signal IO_3_0_IN_pin_0  : std_ulogic := '0';
	signal IO_3_0_IN_pin_1  : std_ulogic := '0';
	signal IO_3_7_IN_pin_0  : std_ulogic := '0';
	signal IO_3_7_IN_pin_1  : std_ulogic := '0';
	signal IO_4_0_IN_pin_0  : std_ulogic := '0';
	signal IO_4_0_IN_pin_1  : std_ulogic := '0';
	signal IO_4_7_IN_pin_0  : std_ulogic := '0';
	signal IO_4_7_IN_pin_1  : std_ulogic := '0';
	signal IO_5_0_IN_pin_0  : std_ulogic := '0';
	signal IO_5_0_IN_pin_1  : std_ulogic := '0';
	signal IO_5_7_IN_pin_0  : std_ulogic := '0';
	signal IO_5_7_IN_pin_1  : std_ulogic := '0';
	signal IO_6_0_IN_pin_0  : std_ulogic := '0';
	signal IO_6_0_IN_pin_1  : std_ulogic := '0';
	signal IO_6_7_IN_pin_0  : std_ulogic := '0';
	signal IO_6_7_IN_pin_1  : std_ulogic := '0';
	signal IO_7_0_IN_pin_0  : std_ulogic := '0';
	signal IO_7_0_IN_pin_1  : std_ulogic := '0';
	signal IO_7_7_IN_pin_0  : std_ulogic := '0';
	signal IO_7_7_IN_pin_1  : std_ulogic := '0';
	signal IO_8_0_IN_pin_0  : std_ulogic := '0';
	signal IO_8_0_IN_pin_1  : std_ulogic := '0';
	signal IO_8_7_IN_pin_0  : std_ulogic := '0';
	signal IO_8_7_IN_pin_1  : std_ulogic := '0';
	signal IO_9_1_IN_pin_0  : std_ulogic := '0';
	signal IO_9_1_IN_pin_1  : std_ulogic := '0';
	signal IO_9_2_IN_pin_0  : std_ulogic := '0';
	signal IO_9_2_IN_pin_1  : std_ulogic := '0';
	signal IO_9_3_IN_pin_0  : std_ulogic := '0';
	signal IO_9_3_IN_pin_1  : std_ulogic := '0';
	signal IO_9_4_IN_pin_0  : std_ulogic := '0';
	signal IO_9_4_IN_pin_1  : std_ulogic := '0';
	signal IO_9_5_IN_pin_0  : std_ulogic := '0';
	signal IO_9_5_IN_pin_1  : std_ulogic := '0';
	signal IO_9_6_IN_pin_0  : std_ulogic := '0';
	signal IO_9_6_IN_pin_1  : std_ulogic := '0';

	-- Tracks --
	signal track_0_1_chanY_n0  : std_ulogic := '0';
	signal track_0_1_chanY_n1  : std_ulogic := '0';
	signal track_0_1_chanY_n10 : std_ulogic := '0';
	signal track_0_1_chanY_n11 : std_ulogic := '0';
	signal track_0_1_chanY_n12 : std_ulogic := '0';
	signal track_0_1_chanY_n13 : std_ulogic := '0';
	signal track_0_1_chanY_n14 : std_ulogic := '0';
	signal track_0_1_chanY_n15 : std_ulogic := '0';
	signal track_0_1_chanY_n2  : std_ulogic := '0';
	signal track_0_1_chanY_n3  : std_ulogic := '0';
	signal track_0_1_chanY_n4  : std_ulogic := '0';
	signal track_0_1_chanY_n5  : std_ulogic := '0';
	signal track_0_1_chanY_n6  : std_ulogic := '0';
	signal track_0_1_chanY_n7  : std_ulogic := '0';
	signal track_0_1_chanY_n8  : std_ulogic := '0';
	signal track_0_1_chanY_n9  : std_ulogic := '0';
	signal track_0_2_chanY_n0  : std_ulogic := '0';
	signal track_0_2_chanY_n1  : std_ulogic := '0';
	signal track_0_2_chanY_n10 : std_ulogic := '0';
	signal track_0_2_chanY_n11 : std_ulogic := '0';
	signal track_0_2_chanY_n12 : std_ulogic := '0';
	signal track_0_2_chanY_n13 : std_ulogic := '0';
	signal track_0_2_chanY_n14 : std_ulogic := '0';
	signal track_0_2_chanY_n15 : std_ulogic := '0';
	signal track_0_2_chanY_n2  : std_ulogic := '0';
	signal track_0_2_chanY_n3  : std_ulogic := '0';
	signal track_0_2_chanY_n4  : std_ulogic := '0';
	signal track_0_2_chanY_n5  : std_ulogic := '0';
	signal track_0_2_chanY_n6  : std_ulogic := '0';
	signal track_0_2_chanY_n7  : std_ulogic := '0';
	signal track_0_2_chanY_n8  : std_ulogic := '0';
	signal track_0_2_chanY_n9  : std_ulogic := '0';
	signal track_0_3_chanY_n0  : std_ulogic := '0';
	signal track_0_3_chanY_n1  : std_ulogic := '0';
	signal track_0_3_chanY_n10 : std_ulogic := '0';
	signal track_0_3_chanY_n11 : std_ulogic := '0';
	signal track_0_3_chanY_n12 : std_ulogic := '0';
	signal track_0_3_chanY_n13 : std_ulogic := '0';
	signal track_0_3_chanY_n14 : std_ulogic := '0';
	signal track_0_3_chanY_n15 : std_ulogic := '0';
	signal track_0_3_chanY_n2  : std_ulogic := '0';
	signal track_0_3_chanY_n3  : std_ulogic := '0';
	signal track_0_3_chanY_n4  : std_ulogic := '0';
	signal track_0_3_chanY_n5  : std_ulogic := '0';
	signal track_0_3_chanY_n6  : std_ulogic := '0';
	signal track_0_3_chanY_n7  : std_ulogic := '0';
	signal track_0_3_chanY_n8  : std_ulogic := '0';
	signal track_0_3_chanY_n9  : std_ulogic := '0';
	signal track_0_4_chanY_n0  : std_ulogic := '0';
	signal track_0_4_chanY_n1  : std_ulogic := '0';
	signal track_0_4_chanY_n10 : std_ulogic := '0';
	signal track_0_4_chanY_n11 : std_ulogic := '0';
	signal track_0_4_chanY_n12 : std_ulogic := '0';
	signal track_0_4_chanY_n13 : std_ulogic := '0';
	signal track_0_4_chanY_n14 : std_ulogic := '0';
	signal track_0_4_chanY_n15 : std_ulogic := '0';
	signal track_0_4_chanY_n2  : std_ulogic := '0';
	signal track_0_4_chanY_n3  : std_ulogic := '0';
	signal track_0_4_chanY_n4  : std_ulogic := '0';
	signal track_0_4_chanY_n5  : std_ulogic := '0';
	signal track_0_4_chanY_n6  : std_ulogic := '0';
	signal track_0_4_chanY_n7  : std_ulogic := '0';
	signal track_0_4_chanY_n8  : std_ulogic := '0';
	signal track_0_4_chanY_n9  : std_ulogic := '0';
	signal track_0_5_chanY_n0  : std_ulogic := '0';
	signal track_0_5_chanY_n1  : std_ulogic := '0';
	signal track_0_5_chanY_n10 : std_ulogic := '0';
	signal track_0_5_chanY_n11 : std_ulogic := '0';
	signal track_0_5_chanY_n12 : std_ulogic := '0';
	signal track_0_5_chanY_n13 : std_ulogic := '0';
	signal track_0_5_chanY_n14 : std_ulogic := '0';
	signal track_0_5_chanY_n15 : std_ulogic := '0';
	signal track_0_5_chanY_n2  : std_ulogic := '0';
	signal track_0_5_chanY_n3  : std_ulogic := '0';
	signal track_0_5_chanY_n4  : std_ulogic := '0';
	signal track_0_5_chanY_n5  : std_ulogic := '0';
	signal track_0_5_chanY_n6  : std_ulogic := '0';
	signal track_0_5_chanY_n7  : std_ulogic := '0';
	signal track_0_5_chanY_n8  : std_ulogic := '0';
	signal track_0_5_chanY_n9  : std_ulogic := '0';
	signal track_0_6_chanY_n0  : std_ulogic := '0';
	signal track_0_6_chanY_n1  : std_ulogic := '0';
	signal track_0_6_chanY_n10 : std_ulogic := '0';
	signal track_0_6_chanY_n11 : std_ulogic := '0';
	signal track_0_6_chanY_n12 : std_ulogic := '0';
	signal track_0_6_chanY_n13 : std_ulogic := '0';
	signal track_0_6_chanY_n14 : std_ulogic := '0';
	signal track_0_6_chanY_n15 : std_ulogic := '0';
	signal track_0_6_chanY_n2  : std_ulogic := '0';
	signal track_0_6_chanY_n3  : std_ulogic := '0';
	signal track_0_6_chanY_n4  : std_ulogic := '0';
	signal track_0_6_chanY_n5  : std_ulogic := '0';
	signal track_0_6_chanY_n6  : std_ulogic := '0';
	signal track_0_6_chanY_n7  : std_ulogic := '0';
	signal track_0_6_chanY_n8  : std_ulogic := '0';
	signal track_0_6_chanY_n9  : std_ulogic := '0';
	signal track_1_0_chanX_n0  : std_ulogic := '0';
	signal track_1_0_chanX_n1  : std_ulogic := '0';
	signal track_1_0_chanX_n10 : std_ulogic := '0';
	signal track_1_0_chanX_n11 : std_ulogic := '0';
	signal track_1_0_chanX_n12 : std_ulogic := '0';
	signal track_1_0_chanX_n13 : std_ulogic := '0';
	signal track_1_0_chanX_n14 : std_ulogic := '0';
	signal track_1_0_chanX_n15 : std_ulogic := '0';
	signal track_1_0_chanX_n2  : std_ulogic := '0';
	signal track_1_0_chanX_n3  : std_ulogic := '0';
	signal track_1_0_chanX_n4  : std_ulogic := '0';
	signal track_1_0_chanX_n5  : std_ulogic := '0';
	signal track_1_0_chanX_n6  : std_ulogic := '0';
	signal track_1_0_chanX_n7  : std_ulogic := '0';
	signal track_1_0_chanX_n8  : std_ulogic := '0';
	signal track_1_0_chanX_n9  : std_ulogic := '0';
	signal track_1_1_chanX_n0  : std_ulogic := '0';
	signal track_1_1_chanX_n1  : std_ulogic := '0';
	signal track_1_1_chanX_n10 : std_ulogic := '0';
	signal track_1_1_chanX_n11 : std_ulogic := '0';
	signal track_1_1_chanX_n12 : std_ulogic := '0';
	signal track_1_1_chanX_n13 : std_ulogic := '0';
	signal track_1_1_chanX_n14 : std_ulogic := '0';
	signal track_1_1_chanX_n15 : std_ulogic := '0';
	signal track_1_1_chanX_n2  : std_ulogic := '0';
	signal track_1_1_chanX_n3  : std_ulogic := '0';
	signal track_1_1_chanX_n4  : std_ulogic := '0';
	signal track_1_1_chanX_n5  : std_ulogic := '0';
	signal track_1_1_chanX_n6  : std_ulogic := '0';
	signal track_1_1_chanX_n7  : std_ulogic := '0';
	signal track_1_1_chanX_n8  : std_ulogic := '0';
	signal track_1_1_chanX_n9  : std_ulogic := '0';
	signal track_1_1_chanY_n0  : std_ulogic := '0';
	signal track_1_1_chanY_n1  : std_ulogic := '0';
	signal track_1_1_chanY_n10 : std_ulogic := '0';
	signal track_1_1_chanY_n11 : std_ulogic := '0';
	signal track_1_1_chanY_n12 : std_ulogic := '0';
	signal track_1_1_chanY_n13 : std_ulogic := '0';
	signal track_1_1_chanY_n14 : std_ulogic := '0';
	signal track_1_1_chanY_n15 : std_ulogic := '0';
	signal track_1_1_chanY_n2  : std_ulogic := '0';
	signal track_1_1_chanY_n3  : std_ulogic := '0';
	signal track_1_1_chanY_n4  : std_ulogic := '0';
	signal track_1_1_chanY_n5  : std_ulogic := '0';
	signal track_1_1_chanY_n6  : std_ulogic := '0';
	signal track_1_1_chanY_n7  : std_ulogic := '0';
	signal track_1_1_chanY_n8  : std_ulogic := '0';
	signal track_1_1_chanY_n9  : std_ulogic := '0';
	signal track_1_2_chanX_n0  : std_ulogic := '0';
	signal track_1_2_chanX_n1  : std_ulogic := '0';
	signal track_1_2_chanX_n10 : std_ulogic := '0';
	signal track_1_2_chanX_n11 : std_ulogic := '0';
	signal track_1_2_chanX_n12 : std_ulogic := '0';
	signal track_1_2_chanX_n13 : std_ulogic := '0';
	signal track_1_2_chanX_n14 : std_ulogic := '0';
	signal track_1_2_chanX_n15 : std_ulogic := '0';
	signal track_1_2_chanX_n2  : std_ulogic := '0';
	signal track_1_2_chanX_n3  : std_ulogic := '0';
	signal track_1_2_chanX_n4  : std_ulogic := '0';
	signal track_1_2_chanX_n5  : std_ulogic := '0';
	signal track_1_2_chanX_n6  : std_ulogic := '0';
	signal track_1_2_chanX_n7  : std_ulogic := '0';
	signal track_1_2_chanX_n8  : std_ulogic := '0';
	signal track_1_2_chanX_n9  : std_ulogic := '0';
	signal track_1_2_chanY_n0  : std_ulogic := '0';
	signal track_1_2_chanY_n1  : std_ulogic := '0';
	signal track_1_2_chanY_n10 : std_ulogic := '0';
	signal track_1_2_chanY_n11 : std_ulogic := '0';
	signal track_1_2_chanY_n12 : std_ulogic := '0';
	signal track_1_2_chanY_n13 : std_ulogic := '0';
	signal track_1_2_chanY_n14 : std_ulogic := '0';
	signal track_1_2_chanY_n15 : std_ulogic := '0';
	signal track_1_2_chanY_n2  : std_ulogic := '0';
	signal track_1_2_chanY_n3  : std_ulogic := '0';
	signal track_1_2_chanY_n4  : std_ulogic := '0';
	signal track_1_2_chanY_n5  : std_ulogic := '0';
	signal track_1_2_chanY_n6  : std_ulogic := '0';
	signal track_1_2_chanY_n7  : std_ulogic := '0';
	signal track_1_2_chanY_n8  : std_ulogic := '0';
	signal track_1_2_chanY_n9  : std_ulogic := '0';
	signal track_1_3_chanX_n0  : std_ulogic := '0';
	signal track_1_3_chanX_n1  : std_ulogic := '0';
	signal track_1_3_chanX_n10 : std_ulogic := '0';
	signal track_1_3_chanX_n11 : std_ulogic := '0';
	signal track_1_3_chanX_n12 : std_ulogic := '0';
	signal track_1_3_chanX_n13 : std_ulogic := '0';
	signal track_1_3_chanX_n14 : std_ulogic := '0';
	signal track_1_3_chanX_n15 : std_ulogic := '0';
	signal track_1_3_chanX_n2  : std_ulogic := '0';
	signal track_1_3_chanX_n3  : std_ulogic := '0';
	signal track_1_3_chanX_n4  : std_ulogic := '0';
	signal track_1_3_chanX_n5  : std_ulogic := '0';
	signal track_1_3_chanX_n6  : std_ulogic := '0';
	signal track_1_3_chanX_n7  : std_ulogic := '0';
	signal track_1_3_chanX_n8  : std_ulogic := '0';
	signal track_1_3_chanX_n9  : std_ulogic := '0';
	signal track_1_3_chanY_n0  : std_ulogic := '0';
	signal track_1_3_chanY_n1  : std_ulogic := '0';
	signal track_1_3_chanY_n10 : std_ulogic := '0';
	signal track_1_3_chanY_n11 : std_ulogic := '0';
	signal track_1_3_chanY_n12 : std_ulogic := '0';
	signal track_1_3_chanY_n13 : std_ulogic := '0';
	signal track_1_3_chanY_n14 : std_ulogic := '0';
	signal track_1_3_chanY_n15 : std_ulogic := '0';
	signal track_1_3_chanY_n2  : std_ulogic := '0';
	signal track_1_3_chanY_n3  : std_ulogic := '0';
	signal track_1_3_chanY_n4  : std_ulogic := '0';
	signal track_1_3_chanY_n5  : std_ulogic := '0';
	signal track_1_3_chanY_n6  : std_ulogic := '0';
	signal track_1_3_chanY_n7  : std_ulogic := '0';
	signal track_1_3_chanY_n8  : std_ulogic := '0';
	signal track_1_3_chanY_n9  : std_ulogic := '0';
	signal track_1_4_chanX_n0  : std_ulogic := '0';
	signal track_1_4_chanX_n1  : std_ulogic := '0';
	signal track_1_4_chanX_n10 : std_ulogic := '0';
	signal track_1_4_chanX_n11 : std_ulogic := '0';
	signal track_1_4_chanX_n12 : std_ulogic := '0';
	signal track_1_4_chanX_n13 : std_ulogic := '0';
	signal track_1_4_chanX_n14 : std_ulogic := '0';
	signal track_1_4_chanX_n15 : std_ulogic := '0';
	signal track_1_4_chanX_n2  : std_ulogic := '0';
	signal track_1_4_chanX_n3  : std_ulogic := '0';
	signal track_1_4_chanX_n4  : std_ulogic := '0';
	signal track_1_4_chanX_n5  : std_ulogic := '0';
	signal track_1_4_chanX_n6  : std_ulogic := '0';
	signal track_1_4_chanX_n7  : std_ulogic := '0';
	signal track_1_4_chanX_n8  : std_ulogic := '0';
	signal track_1_4_chanX_n9  : std_ulogic := '0';
	signal track_1_4_chanY_n0  : std_ulogic := '0';
	signal track_1_4_chanY_n1  : std_ulogic := '0';
	signal track_1_4_chanY_n10 : std_ulogic := '0';
	signal track_1_4_chanY_n11 : std_ulogic := '0';
	signal track_1_4_chanY_n12 : std_ulogic := '0';
	signal track_1_4_chanY_n13 : std_ulogic := '0';
	signal track_1_4_chanY_n14 : std_ulogic := '0';
	signal track_1_4_chanY_n15 : std_ulogic := '0';
	signal track_1_4_chanY_n2  : std_ulogic := '0';
	signal track_1_4_chanY_n3  : std_ulogic := '0';
	signal track_1_4_chanY_n4  : std_ulogic := '0';
	signal track_1_4_chanY_n5  : std_ulogic := '0';
	signal track_1_4_chanY_n6  : std_ulogic := '0';
	signal track_1_4_chanY_n7  : std_ulogic := '0';
	signal track_1_4_chanY_n8  : std_ulogic := '0';
	signal track_1_4_chanY_n9  : std_ulogic := '0';
	signal track_1_5_chanX_n0  : std_ulogic := '0';
	signal track_1_5_chanX_n1  : std_ulogic := '0';
	signal track_1_5_chanX_n10 : std_ulogic := '0';
	signal track_1_5_chanX_n11 : std_ulogic := '0';
	signal track_1_5_chanX_n12 : std_ulogic := '0';
	signal track_1_5_chanX_n13 : std_ulogic := '0';
	signal track_1_5_chanX_n14 : std_ulogic := '0';
	signal track_1_5_chanX_n15 : std_ulogic := '0';
	signal track_1_5_chanX_n2  : std_ulogic := '0';
	signal track_1_5_chanX_n3  : std_ulogic := '0';
	signal track_1_5_chanX_n4  : std_ulogic := '0';
	signal track_1_5_chanX_n5  : std_ulogic := '0';
	signal track_1_5_chanX_n6  : std_ulogic := '0';
	signal track_1_5_chanX_n7  : std_ulogic := '0';
	signal track_1_5_chanX_n8  : std_ulogic := '0';
	signal track_1_5_chanX_n9  : std_ulogic := '0';
	signal track_1_5_chanY_n0  : std_ulogic := '0';
	signal track_1_5_chanY_n1  : std_ulogic := '0';
	signal track_1_5_chanY_n10 : std_ulogic := '0';
	signal track_1_5_chanY_n11 : std_ulogic := '0';
	signal track_1_5_chanY_n12 : std_ulogic := '0';
	signal track_1_5_chanY_n13 : std_ulogic := '0';
	signal track_1_5_chanY_n14 : std_ulogic := '0';
	signal track_1_5_chanY_n15 : std_ulogic := '0';
	signal track_1_5_chanY_n2  : std_ulogic := '0';
	signal track_1_5_chanY_n3  : std_ulogic := '0';
	signal track_1_5_chanY_n4  : std_ulogic := '0';
	signal track_1_5_chanY_n5  : std_ulogic := '0';
	signal track_1_5_chanY_n6  : std_ulogic := '0';
	signal track_1_5_chanY_n7  : std_ulogic := '0';
	signal track_1_5_chanY_n8  : std_ulogic := '0';
	signal track_1_5_chanY_n9  : std_ulogic := '0';
	signal track_1_6_chanX_n0  : std_ulogic := '0';
	signal track_1_6_chanX_n1  : std_ulogic := '0';
	signal track_1_6_chanX_n10 : std_ulogic := '0';
	signal track_1_6_chanX_n11 : std_ulogic := '0';
	signal track_1_6_chanX_n12 : std_ulogic := '0';
	signal track_1_6_chanX_n13 : std_ulogic := '0';
	signal track_1_6_chanX_n14 : std_ulogic := '0';
	signal track_1_6_chanX_n15 : std_ulogic := '0';
	signal track_1_6_chanX_n2  : std_ulogic := '0';
	signal track_1_6_chanX_n3  : std_ulogic := '0';
	signal track_1_6_chanX_n4  : std_ulogic := '0';
	signal track_1_6_chanX_n5  : std_ulogic := '0';
	signal track_1_6_chanX_n6  : std_ulogic := '0';
	signal track_1_6_chanX_n7  : std_ulogic := '0';
	signal track_1_6_chanX_n8  : std_ulogic := '0';
	signal track_1_6_chanX_n9  : std_ulogic := '0';
	signal track_1_6_chanY_n0  : std_ulogic := '0';
	signal track_1_6_chanY_n1  : std_ulogic := '0';
	signal track_1_6_chanY_n10 : std_ulogic := '0';
	signal track_1_6_chanY_n11 : std_ulogic := '0';
	signal track_1_6_chanY_n12 : std_ulogic := '0';
	signal track_1_6_chanY_n13 : std_ulogic := '0';
	signal track_1_6_chanY_n14 : std_ulogic := '0';
	signal track_1_6_chanY_n15 : std_ulogic := '0';
	signal track_1_6_chanY_n2  : std_ulogic := '0';
	signal track_1_6_chanY_n3  : std_ulogic := '0';
	signal track_1_6_chanY_n4  : std_ulogic := '0';
	signal track_1_6_chanY_n5  : std_ulogic := '0';
	signal track_1_6_chanY_n6  : std_ulogic := '0';
	signal track_1_6_chanY_n7  : std_ulogic := '0';
	signal track_1_6_chanY_n8  : std_ulogic := '0';
	signal track_1_6_chanY_n9  : std_ulogic := '0';
	signal track_2_0_chanX_n0  : std_ulogic := '0';
	signal track_2_0_chanX_n1  : std_ulogic := '0';
	signal track_2_0_chanX_n10 : std_ulogic := '0';
	signal track_2_0_chanX_n11 : std_ulogic := '0';
	signal track_2_0_chanX_n12 : std_ulogic := '0';
	signal track_2_0_chanX_n13 : std_ulogic := '0';
	signal track_2_0_chanX_n14 : std_ulogic := '0';
	signal track_2_0_chanX_n15 : std_ulogic := '0';
	signal track_2_0_chanX_n2  : std_ulogic := '0';
	signal track_2_0_chanX_n3  : std_ulogic := '0';
	signal track_2_0_chanX_n4  : std_ulogic := '0';
	signal track_2_0_chanX_n5  : std_ulogic := '0';
	signal track_2_0_chanX_n6  : std_ulogic := '0';
	signal track_2_0_chanX_n7  : std_ulogic := '0';
	signal track_2_0_chanX_n8  : std_ulogic := '0';
	signal track_2_0_chanX_n9  : std_ulogic := '0';
	signal track_2_1_chanX_n0  : std_ulogic := '0';
	signal track_2_1_chanX_n1  : std_ulogic := '0';
	signal track_2_1_chanX_n10 : std_ulogic := '0';
	signal track_2_1_chanX_n11 : std_ulogic := '0';
	signal track_2_1_chanX_n12 : std_ulogic := '0';
	signal track_2_1_chanX_n13 : std_ulogic := '0';
	signal track_2_1_chanX_n14 : std_ulogic := '0';
	signal track_2_1_chanX_n15 : std_ulogic := '0';
	signal track_2_1_chanX_n2  : std_ulogic := '0';
	signal track_2_1_chanX_n3  : std_ulogic := '0';
	signal track_2_1_chanX_n4  : std_ulogic := '0';
	signal track_2_1_chanX_n5  : std_ulogic := '0';
	signal track_2_1_chanX_n6  : std_ulogic := '0';
	signal track_2_1_chanX_n7  : std_ulogic := '0';
	signal track_2_1_chanX_n8  : std_ulogic := '0';
	signal track_2_1_chanX_n9  : std_ulogic := '0';
	signal track_2_1_chanY_n0  : std_ulogic := '0';
	signal track_2_1_chanY_n1  : std_ulogic := '0';
	signal track_2_1_chanY_n10 : std_ulogic := '0';
	signal track_2_1_chanY_n11 : std_ulogic := '0';
	signal track_2_1_chanY_n12 : std_ulogic := '0';
	signal track_2_1_chanY_n13 : std_ulogic := '0';
	signal track_2_1_chanY_n14 : std_ulogic := '0';
	signal track_2_1_chanY_n15 : std_ulogic := '0';
	signal track_2_1_chanY_n2  : std_ulogic := '0';
	signal track_2_1_chanY_n3  : std_ulogic := '0';
	signal track_2_1_chanY_n4  : std_ulogic := '0';
	signal track_2_1_chanY_n5  : std_ulogic := '0';
	signal track_2_1_chanY_n6  : std_ulogic := '0';
	signal track_2_1_chanY_n7  : std_ulogic := '0';
	signal track_2_1_chanY_n8  : std_ulogic := '0';
	signal track_2_1_chanY_n9  : std_ulogic := '0';
	signal track_2_2_chanX_n0  : std_ulogic := '0';
	signal track_2_2_chanX_n1  : std_ulogic := '0';
	signal track_2_2_chanX_n10 : std_ulogic := '0';
	signal track_2_2_chanX_n11 : std_ulogic := '0';
	signal track_2_2_chanX_n12 : std_ulogic := '0';
	signal track_2_2_chanX_n13 : std_ulogic := '0';
	signal track_2_2_chanX_n14 : std_ulogic := '0';
	signal track_2_2_chanX_n15 : std_ulogic := '0';
	signal track_2_2_chanX_n2  : std_ulogic := '0';
	signal track_2_2_chanX_n3  : std_ulogic := '0';
	signal track_2_2_chanX_n4  : std_ulogic := '0';
	signal track_2_2_chanX_n5  : std_ulogic := '0';
	signal track_2_2_chanX_n6  : std_ulogic := '0';
	signal track_2_2_chanX_n7  : std_ulogic := '0';
	signal track_2_2_chanX_n8  : std_ulogic := '0';
	signal track_2_2_chanX_n9  : std_ulogic := '0';
	signal track_2_2_chanY_n0  : std_ulogic := '0';
	signal track_2_2_chanY_n1  : std_ulogic := '0';
	signal track_2_2_chanY_n10 : std_ulogic := '0';
	signal track_2_2_chanY_n11 : std_ulogic := '0';
	signal track_2_2_chanY_n12 : std_ulogic := '0';
	signal track_2_2_chanY_n13 : std_ulogic := '0';
	signal track_2_2_chanY_n14 : std_ulogic := '0';
	signal track_2_2_chanY_n15 : std_ulogic := '0';
	signal track_2_2_chanY_n2  : std_ulogic := '0';
	signal track_2_2_chanY_n3  : std_ulogic := '0';
	signal track_2_2_chanY_n4  : std_ulogic := '0';
	signal track_2_2_chanY_n5  : std_ulogic := '0';
	signal track_2_2_chanY_n6  : std_ulogic := '0';
	signal track_2_2_chanY_n7  : std_ulogic := '0';
	signal track_2_2_chanY_n8  : std_ulogic := '0';
	signal track_2_2_chanY_n9  : std_ulogic := '0';
	signal track_2_3_chanX_n0  : std_ulogic := '0';
	signal track_2_3_chanX_n1  : std_ulogic := '0';
	signal track_2_3_chanX_n10 : std_ulogic := '0';
	signal track_2_3_chanX_n11 : std_ulogic := '0';
	signal track_2_3_chanX_n12 : std_ulogic := '0';
	signal track_2_3_chanX_n13 : std_ulogic := '0';
	signal track_2_3_chanX_n14 : std_ulogic := '0';
	signal track_2_3_chanX_n15 : std_ulogic := '0';
	signal track_2_3_chanX_n2  : std_ulogic := '0';
	signal track_2_3_chanX_n3  : std_ulogic := '0';
	signal track_2_3_chanX_n4  : std_ulogic := '0';
	signal track_2_3_chanX_n5  : std_ulogic := '0';
	signal track_2_3_chanX_n6  : std_ulogic := '0';
	signal track_2_3_chanX_n7  : std_ulogic := '0';
	signal track_2_3_chanX_n8  : std_ulogic := '0';
	signal track_2_3_chanX_n9  : std_ulogic := '0';
	signal track_2_3_chanY_n0  : std_ulogic := '0';
	signal track_2_3_chanY_n1  : std_ulogic := '0';
	signal track_2_3_chanY_n10 : std_ulogic := '0';
	signal track_2_3_chanY_n11 : std_ulogic := '0';
	signal track_2_3_chanY_n12 : std_ulogic := '0';
	signal track_2_3_chanY_n13 : std_ulogic := '0';
	signal track_2_3_chanY_n14 : std_ulogic := '0';
	signal track_2_3_chanY_n15 : std_ulogic := '0';
	signal track_2_3_chanY_n2  : std_ulogic := '0';
	signal track_2_3_chanY_n3  : std_ulogic := '0';
	signal track_2_3_chanY_n4  : std_ulogic := '0';
	signal track_2_3_chanY_n5  : std_ulogic := '0';
	signal track_2_3_chanY_n6  : std_ulogic := '0';
	signal track_2_3_chanY_n7  : std_ulogic := '0';
	signal track_2_3_chanY_n8  : std_ulogic := '0';
	signal track_2_3_chanY_n9  : std_ulogic := '0';
	signal track_2_4_chanX_n0  : std_ulogic := '0';
	signal track_2_4_chanX_n1  : std_ulogic := '0';
	signal track_2_4_chanX_n10 : std_ulogic := '0';
	signal track_2_4_chanX_n11 : std_ulogic := '0';
	signal track_2_4_chanX_n12 : std_ulogic := '0';
	signal track_2_4_chanX_n13 : std_ulogic := '0';
	signal track_2_4_chanX_n14 : std_ulogic := '0';
	signal track_2_4_chanX_n15 : std_ulogic := '0';
	signal track_2_4_chanX_n2  : std_ulogic := '0';
	signal track_2_4_chanX_n3  : std_ulogic := '0';
	signal track_2_4_chanX_n4  : std_ulogic := '0';
	signal track_2_4_chanX_n5  : std_ulogic := '0';
	signal track_2_4_chanX_n6  : std_ulogic := '0';
	signal track_2_4_chanX_n7  : std_ulogic := '0';
	signal track_2_4_chanX_n8  : std_ulogic := '0';
	signal track_2_4_chanX_n9  : std_ulogic := '0';
	signal track_2_4_chanY_n0  : std_ulogic := '0';
	signal track_2_4_chanY_n1  : std_ulogic := '0';
	signal track_2_4_chanY_n10 : std_ulogic := '0';
	signal track_2_4_chanY_n11 : std_ulogic := '0';
	signal track_2_4_chanY_n12 : std_ulogic := '0';
	signal track_2_4_chanY_n13 : std_ulogic := '0';
	signal track_2_4_chanY_n14 : std_ulogic := '0';
	signal track_2_4_chanY_n15 : std_ulogic := '0';
	signal track_2_4_chanY_n2  : std_ulogic := '0';
	signal track_2_4_chanY_n3  : std_ulogic := '0';
	signal track_2_4_chanY_n4  : std_ulogic := '0';
	signal track_2_4_chanY_n5  : std_ulogic := '0';
	signal track_2_4_chanY_n6  : std_ulogic := '0';
	signal track_2_4_chanY_n7  : std_ulogic := '0';
	signal track_2_4_chanY_n8  : std_ulogic := '0';
	signal track_2_4_chanY_n9  : std_ulogic := '0';
	signal track_2_5_chanX_n0  : std_ulogic := '0';
	signal track_2_5_chanX_n1  : std_ulogic := '0';
	signal track_2_5_chanX_n10 : std_ulogic := '0';
	signal track_2_5_chanX_n11 : std_ulogic := '0';
	signal track_2_5_chanX_n12 : std_ulogic := '0';
	signal track_2_5_chanX_n13 : std_ulogic := '0';
	signal track_2_5_chanX_n14 : std_ulogic := '0';
	signal track_2_5_chanX_n15 : std_ulogic := '0';
	signal track_2_5_chanX_n2  : std_ulogic := '0';
	signal track_2_5_chanX_n3  : std_ulogic := '0';
	signal track_2_5_chanX_n4  : std_ulogic := '0';
	signal track_2_5_chanX_n5  : std_ulogic := '0';
	signal track_2_5_chanX_n6  : std_ulogic := '0';
	signal track_2_5_chanX_n7  : std_ulogic := '0';
	signal track_2_5_chanX_n8  : std_ulogic := '0';
	signal track_2_5_chanX_n9  : std_ulogic := '0';
	signal track_2_5_chanY_n0  : std_ulogic := '0';
	signal track_2_5_chanY_n1  : std_ulogic := '0';
	signal track_2_5_chanY_n10 : std_ulogic := '0';
	signal track_2_5_chanY_n11 : std_ulogic := '0';
	signal track_2_5_chanY_n12 : std_ulogic := '0';
	signal track_2_5_chanY_n13 : std_ulogic := '0';
	signal track_2_5_chanY_n14 : std_ulogic := '0';
	signal track_2_5_chanY_n15 : std_ulogic := '0';
	signal track_2_5_chanY_n2  : std_ulogic := '0';
	signal track_2_5_chanY_n3  : std_ulogic := '0';
	signal track_2_5_chanY_n4  : std_ulogic := '0';
	signal track_2_5_chanY_n5  : std_ulogic := '0';
	signal track_2_5_chanY_n6  : std_ulogic := '0';
	signal track_2_5_chanY_n7  : std_ulogic := '0';
	signal track_2_5_chanY_n8  : std_ulogic := '0';
	signal track_2_5_chanY_n9  : std_ulogic := '0';
	signal track_2_6_chanX_n0  : std_ulogic := '0';
	signal track_2_6_chanX_n1  : std_ulogic := '0';
	signal track_2_6_chanX_n10 : std_ulogic := '0';
	signal track_2_6_chanX_n11 : std_ulogic := '0';
	signal track_2_6_chanX_n12 : std_ulogic := '0';
	signal track_2_6_chanX_n13 : std_ulogic := '0';
	signal track_2_6_chanX_n14 : std_ulogic := '0';
	signal track_2_6_chanX_n15 : std_ulogic := '0';
	signal track_2_6_chanX_n2  : std_ulogic := '0';
	signal track_2_6_chanX_n3  : std_ulogic := '0';
	signal track_2_6_chanX_n4  : std_ulogic := '0';
	signal track_2_6_chanX_n5  : std_ulogic := '0';
	signal track_2_6_chanX_n6  : std_ulogic := '0';
	signal track_2_6_chanX_n7  : std_ulogic := '0';
	signal track_2_6_chanX_n8  : std_ulogic := '0';
	signal track_2_6_chanX_n9  : std_ulogic := '0';
	signal track_2_6_chanY_n0  : std_ulogic := '0';
	signal track_2_6_chanY_n1  : std_ulogic := '0';
	signal track_2_6_chanY_n10 : std_ulogic := '0';
	signal track_2_6_chanY_n11 : std_ulogic := '0';
	signal track_2_6_chanY_n12 : std_ulogic := '0';
	signal track_2_6_chanY_n13 : std_ulogic := '0';
	signal track_2_6_chanY_n14 : std_ulogic := '0';
	signal track_2_6_chanY_n15 : std_ulogic := '0';
	signal track_2_6_chanY_n2  : std_ulogic := '0';
	signal track_2_6_chanY_n3  : std_ulogic := '0';
	signal track_2_6_chanY_n4  : std_ulogic := '0';
	signal track_2_6_chanY_n5  : std_ulogic := '0';
	signal track_2_6_chanY_n6  : std_ulogic := '0';
	signal track_2_6_chanY_n7  : std_ulogic := '0';
	signal track_2_6_chanY_n8  : std_ulogic := '0';
	signal track_2_6_chanY_n9  : std_ulogic := '0';
	signal track_3_0_chanX_n0  : std_ulogic := '0';
	signal track_3_0_chanX_n1  : std_ulogic := '0';
	signal track_3_0_chanX_n10 : std_ulogic := '0';
	signal track_3_0_chanX_n11 : std_ulogic := '0';
	signal track_3_0_chanX_n12 : std_ulogic := '0';
	signal track_3_0_chanX_n13 : std_ulogic := '0';
	signal track_3_0_chanX_n14 : std_ulogic := '0';
	signal track_3_0_chanX_n15 : std_ulogic := '0';
	signal track_3_0_chanX_n2  : std_ulogic := '0';
	signal track_3_0_chanX_n3  : std_ulogic := '0';
	signal track_3_0_chanX_n4  : std_ulogic := '0';
	signal track_3_0_chanX_n5  : std_ulogic := '0';
	signal track_3_0_chanX_n6  : std_ulogic := '0';
	signal track_3_0_chanX_n7  : std_ulogic := '0';
	signal track_3_0_chanX_n8  : std_ulogic := '0';
	signal track_3_0_chanX_n9  : std_ulogic := '0';
	signal track_3_1_chanX_n0  : std_ulogic := '0';
	signal track_3_1_chanX_n1  : std_ulogic := '0';
	signal track_3_1_chanX_n10 : std_ulogic := '0';
	signal track_3_1_chanX_n11 : std_ulogic := '0';
	signal track_3_1_chanX_n12 : std_ulogic := '0';
	signal track_3_1_chanX_n13 : std_ulogic := '0';
	signal track_3_1_chanX_n14 : std_ulogic := '0';
	signal track_3_1_chanX_n15 : std_ulogic := '0';
	signal track_3_1_chanX_n2  : std_ulogic := '0';
	signal track_3_1_chanX_n3  : std_ulogic := '0';
	signal track_3_1_chanX_n4  : std_ulogic := '0';
	signal track_3_1_chanX_n5  : std_ulogic := '0';
	signal track_3_1_chanX_n6  : std_ulogic := '0';
	signal track_3_1_chanX_n7  : std_ulogic := '0';
	signal track_3_1_chanX_n8  : std_ulogic := '0';
	signal track_3_1_chanX_n9  : std_ulogic := '0';
	signal track_3_1_chanY_n0  : std_ulogic := '0';
	signal track_3_1_chanY_n1  : std_ulogic := '0';
	signal track_3_1_chanY_n10 : std_ulogic := '0';
	signal track_3_1_chanY_n11 : std_ulogic := '0';
	signal track_3_1_chanY_n12 : std_ulogic := '0';
	signal track_3_1_chanY_n13 : std_ulogic := '0';
	signal track_3_1_chanY_n14 : std_ulogic := '0';
	signal track_3_1_chanY_n15 : std_ulogic := '0';
	signal track_3_1_chanY_n2  : std_ulogic := '0';
	signal track_3_1_chanY_n3  : std_ulogic := '0';
	signal track_3_1_chanY_n4  : std_ulogic := '0';
	signal track_3_1_chanY_n5  : std_ulogic := '0';
	signal track_3_1_chanY_n6  : std_ulogic := '0';
	signal track_3_1_chanY_n7  : std_ulogic := '0';
	signal track_3_1_chanY_n8  : std_ulogic := '0';
	signal track_3_1_chanY_n9  : std_ulogic := '0';
	signal track_3_2_chanX_n0  : std_ulogic := '0';
	signal track_3_2_chanX_n1  : std_ulogic := '0';
	signal track_3_2_chanX_n10 : std_ulogic := '0';
	signal track_3_2_chanX_n11 : std_ulogic := '0';
	signal track_3_2_chanX_n12 : std_ulogic := '0';
	signal track_3_2_chanX_n13 : std_ulogic := '0';
	signal track_3_2_chanX_n14 : std_ulogic := '0';
	signal track_3_2_chanX_n15 : std_ulogic := '0';
	signal track_3_2_chanX_n2  : std_ulogic := '0';
	signal track_3_2_chanX_n3  : std_ulogic := '0';
	signal track_3_2_chanX_n4  : std_ulogic := '0';
	signal track_3_2_chanX_n5  : std_ulogic := '0';
	signal track_3_2_chanX_n6  : std_ulogic := '0';
	signal track_3_2_chanX_n7  : std_ulogic := '0';
	signal track_3_2_chanX_n8  : std_ulogic := '0';
	signal track_3_2_chanX_n9  : std_ulogic := '0';
	signal track_3_2_chanY_n0  : std_ulogic := '0';
	signal track_3_2_chanY_n1  : std_ulogic := '0';
	signal track_3_2_chanY_n10 : std_ulogic := '0';
	signal track_3_2_chanY_n11 : std_ulogic := '0';
	signal track_3_2_chanY_n12 : std_ulogic := '0';
	signal track_3_2_chanY_n13 : std_ulogic := '0';
	signal track_3_2_chanY_n14 : std_ulogic := '0';
	signal track_3_2_chanY_n15 : std_ulogic := '0';
	signal track_3_2_chanY_n2  : std_ulogic := '0';
	signal track_3_2_chanY_n3  : std_ulogic := '0';
	signal track_3_2_chanY_n4  : std_ulogic := '0';
	signal track_3_2_chanY_n5  : std_ulogic := '0';
	signal track_3_2_chanY_n6  : std_ulogic := '0';
	signal track_3_2_chanY_n7  : std_ulogic := '0';
	signal track_3_2_chanY_n8  : std_ulogic := '0';
	signal track_3_2_chanY_n9  : std_ulogic := '0';
	signal track_3_3_chanX_n0  : std_ulogic := '0';
	signal track_3_3_chanX_n1  : std_ulogic := '0';
	signal track_3_3_chanX_n10 : std_ulogic := '0';
	signal track_3_3_chanX_n11 : std_ulogic := '0';
	signal track_3_3_chanX_n12 : std_ulogic := '0';
	signal track_3_3_chanX_n13 : std_ulogic := '0';
	signal track_3_3_chanX_n14 : std_ulogic := '0';
	signal track_3_3_chanX_n15 : std_ulogic := '0';
	signal track_3_3_chanX_n2  : std_ulogic := '0';
	signal track_3_3_chanX_n3  : std_ulogic := '0';
	signal track_3_3_chanX_n4  : std_ulogic := '0';
	signal track_3_3_chanX_n5  : std_ulogic := '0';
	signal track_3_3_chanX_n6  : std_ulogic := '0';
	signal track_3_3_chanX_n7  : std_ulogic := '0';
	signal track_3_3_chanX_n8  : std_ulogic := '0';
	signal track_3_3_chanX_n9  : std_ulogic := '0';
	signal track_3_3_chanY_n0  : std_ulogic := '0';
	signal track_3_3_chanY_n1  : std_ulogic := '0';
	signal track_3_3_chanY_n10 : std_ulogic := '0';
	signal track_3_3_chanY_n11 : std_ulogic := '0';
	signal track_3_3_chanY_n12 : std_ulogic := '0';
	signal track_3_3_chanY_n13 : std_ulogic := '0';
	signal track_3_3_chanY_n14 : std_ulogic := '0';
	signal track_3_3_chanY_n15 : std_ulogic := '0';
	signal track_3_3_chanY_n2  : std_ulogic := '0';
	signal track_3_3_chanY_n3  : std_ulogic := '0';
	signal track_3_3_chanY_n4  : std_ulogic := '0';
	signal track_3_3_chanY_n5  : std_ulogic := '0';
	signal track_3_3_chanY_n6  : std_ulogic := '0';
	signal track_3_3_chanY_n7  : std_ulogic := '0';
	signal track_3_3_chanY_n8  : std_ulogic := '0';
	signal track_3_3_chanY_n9  : std_ulogic := '0';
	signal track_3_4_chanX_n0  : std_ulogic := '0';
	signal track_3_4_chanX_n1  : std_ulogic := '0';
	signal track_3_4_chanX_n10 : std_ulogic := '0';
	signal track_3_4_chanX_n11 : std_ulogic := '0';
	signal track_3_4_chanX_n12 : std_ulogic := '0';
	signal track_3_4_chanX_n13 : std_ulogic := '0';
	signal track_3_4_chanX_n14 : std_ulogic := '0';
	signal track_3_4_chanX_n15 : std_ulogic := '0';
	signal track_3_4_chanX_n2  : std_ulogic := '0';
	signal track_3_4_chanX_n3  : std_ulogic := '0';
	signal track_3_4_chanX_n4  : std_ulogic := '0';
	signal track_3_4_chanX_n5  : std_ulogic := '0';
	signal track_3_4_chanX_n6  : std_ulogic := '0';
	signal track_3_4_chanX_n7  : std_ulogic := '0';
	signal track_3_4_chanX_n8  : std_ulogic := '0';
	signal track_3_4_chanX_n9  : std_ulogic := '0';
	signal track_3_4_chanY_n0  : std_ulogic := '0';
	signal track_3_4_chanY_n1  : std_ulogic := '0';
	signal track_3_4_chanY_n10 : std_ulogic := '0';
	signal track_3_4_chanY_n11 : std_ulogic := '0';
	signal track_3_4_chanY_n12 : std_ulogic := '0';
	signal track_3_4_chanY_n13 : std_ulogic := '0';
	signal track_3_4_chanY_n14 : std_ulogic := '0';
	signal track_3_4_chanY_n15 : std_ulogic := '0';
	signal track_3_4_chanY_n2  : std_ulogic := '0';
	signal track_3_4_chanY_n3  : std_ulogic := '0';
	signal track_3_4_chanY_n4  : std_ulogic := '0';
	signal track_3_4_chanY_n5  : std_ulogic := '0';
	signal track_3_4_chanY_n6  : std_ulogic := '0';
	signal track_3_4_chanY_n7  : std_ulogic := '0';
	signal track_3_4_chanY_n8  : std_ulogic := '0';
	signal track_3_4_chanY_n9  : std_ulogic := '0';
	signal track_3_5_chanX_n0  : std_ulogic := '0';
	signal track_3_5_chanX_n1  : std_ulogic := '0';
	signal track_3_5_chanX_n10 : std_ulogic := '0';
	signal track_3_5_chanX_n11 : std_ulogic := '0';
	signal track_3_5_chanX_n12 : std_ulogic := '0';
	signal track_3_5_chanX_n13 : std_ulogic := '0';
	signal track_3_5_chanX_n14 : std_ulogic := '0';
	signal track_3_5_chanX_n15 : std_ulogic := '0';
	signal track_3_5_chanX_n2  : std_ulogic := '0';
	signal track_3_5_chanX_n3  : std_ulogic := '0';
	signal track_3_5_chanX_n4  : std_ulogic := '0';
	signal track_3_5_chanX_n5  : std_ulogic := '0';
	signal track_3_5_chanX_n6  : std_ulogic := '0';
	signal track_3_5_chanX_n7  : std_ulogic := '0';
	signal track_3_5_chanX_n8  : std_ulogic := '0';
	signal track_3_5_chanX_n9  : std_ulogic := '0';
	signal track_3_5_chanY_n0  : std_ulogic := '0';
	signal track_3_5_chanY_n1  : std_ulogic := '0';
	signal track_3_5_chanY_n10 : std_ulogic := '0';
	signal track_3_5_chanY_n11 : std_ulogic := '0';
	signal track_3_5_chanY_n12 : std_ulogic := '0';
	signal track_3_5_chanY_n13 : std_ulogic := '0';
	signal track_3_5_chanY_n14 : std_ulogic := '0';
	signal track_3_5_chanY_n15 : std_ulogic := '0';
	signal track_3_5_chanY_n2  : std_ulogic := '0';
	signal track_3_5_chanY_n3  : std_ulogic := '0';
	signal track_3_5_chanY_n4  : std_ulogic := '0';
	signal track_3_5_chanY_n5  : std_ulogic := '0';
	signal track_3_5_chanY_n6  : std_ulogic := '0';
	signal track_3_5_chanY_n7  : std_ulogic := '0';
	signal track_3_5_chanY_n8  : std_ulogic := '0';
	signal track_3_5_chanY_n9  : std_ulogic := '0';
	signal track_3_6_chanX_n0  : std_ulogic := '0';
	signal track_3_6_chanX_n1  : std_ulogic := '0';
	signal track_3_6_chanX_n10 : std_ulogic := '0';
	signal track_3_6_chanX_n11 : std_ulogic := '0';
	signal track_3_6_chanX_n12 : std_ulogic := '0';
	signal track_3_6_chanX_n13 : std_ulogic := '0';
	signal track_3_6_chanX_n14 : std_ulogic := '0';
	signal track_3_6_chanX_n15 : std_ulogic := '0';
	signal track_3_6_chanX_n2  : std_ulogic := '0';
	signal track_3_6_chanX_n3  : std_ulogic := '0';
	signal track_3_6_chanX_n4  : std_ulogic := '0';
	signal track_3_6_chanX_n5  : std_ulogic := '0';
	signal track_3_6_chanX_n6  : std_ulogic := '0';
	signal track_3_6_chanX_n7  : std_ulogic := '0';
	signal track_3_6_chanX_n8  : std_ulogic := '0';
	signal track_3_6_chanX_n9  : std_ulogic := '0';
	signal track_3_6_chanY_n0  : std_ulogic := '0';
	signal track_3_6_chanY_n1  : std_ulogic := '0';
	signal track_3_6_chanY_n10 : std_ulogic := '0';
	signal track_3_6_chanY_n11 : std_ulogic := '0';
	signal track_3_6_chanY_n12 : std_ulogic := '0';
	signal track_3_6_chanY_n13 : std_ulogic := '0';
	signal track_3_6_chanY_n14 : std_ulogic := '0';
	signal track_3_6_chanY_n15 : std_ulogic := '0';
	signal track_3_6_chanY_n2  : std_ulogic := '0';
	signal track_3_6_chanY_n3  : std_ulogic := '0';
	signal track_3_6_chanY_n4  : std_ulogic := '0';
	signal track_3_6_chanY_n5  : std_ulogic := '0';
	signal track_3_6_chanY_n6  : std_ulogic := '0';
	signal track_3_6_chanY_n7  : std_ulogic := '0';
	signal track_3_6_chanY_n8  : std_ulogic := '0';
	signal track_3_6_chanY_n9  : std_ulogic := '0';
	signal track_4_0_chanX_n0  : std_ulogic := '0';
	signal track_4_0_chanX_n1  : std_ulogic := '0';
	signal track_4_0_chanX_n10 : std_ulogic := '0';
	signal track_4_0_chanX_n11 : std_ulogic := '0';
	signal track_4_0_chanX_n12 : std_ulogic := '0';
	signal track_4_0_chanX_n13 : std_ulogic := '0';
	signal track_4_0_chanX_n14 : std_ulogic := '0';
	signal track_4_0_chanX_n15 : std_ulogic := '0';
	signal track_4_0_chanX_n2  : std_ulogic := '0';
	signal track_4_0_chanX_n3  : std_ulogic := '0';
	signal track_4_0_chanX_n4  : std_ulogic := '0';
	signal track_4_0_chanX_n5  : std_ulogic := '0';
	signal track_4_0_chanX_n6  : std_ulogic := '0';
	signal track_4_0_chanX_n7  : std_ulogic := '0';
	signal track_4_0_chanX_n8  : std_ulogic := '0';
	signal track_4_0_chanX_n9  : std_ulogic := '0';
	signal track_4_1_chanX_n0  : std_ulogic := '0';
	signal track_4_1_chanX_n1  : std_ulogic := '0';
	signal track_4_1_chanX_n10 : std_ulogic := '0';
	signal track_4_1_chanX_n11 : std_ulogic := '0';
	signal track_4_1_chanX_n12 : std_ulogic := '0';
	signal track_4_1_chanX_n13 : std_ulogic := '0';
	signal track_4_1_chanX_n14 : std_ulogic := '0';
	signal track_4_1_chanX_n15 : std_ulogic := '0';
	signal track_4_1_chanX_n2  : std_ulogic := '0';
	signal track_4_1_chanX_n3  : std_ulogic := '0';
	signal track_4_1_chanX_n4  : std_ulogic := '0';
	signal track_4_1_chanX_n5  : std_ulogic := '0';
	signal track_4_1_chanX_n6  : std_ulogic := '0';
	signal track_4_1_chanX_n7  : std_ulogic := '0';
	signal track_4_1_chanX_n8  : std_ulogic := '0';
	signal track_4_1_chanX_n9  : std_ulogic := '0';
	signal track_4_1_chanY_n0  : std_ulogic := '0';
	signal track_4_1_chanY_n1  : std_ulogic := '0';
	signal track_4_1_chanY_n10 : std_ulogic := '0';
	signal track_4_1_chanY_n11 : std_ulogic := '0';
	signal track_4_1_chanY_n12 : std_ulogic := '0';
	signal track_4_1_chanY_n13 : std_ulogic := '0';
	signal track_4_1_chanY_n14 : std_ulogic := '0';
	signal track_4_1_chanY_n15 : std_ulogic := '0';
	signal track_4_1_chanY_n2  : std_ulogic := '0';
	signal track_4_1_chanY_n3  : std_ulogic := '0';
	signal track_4_1_chanY_n4  : std_ulogic := '0';
	signal track_4_1_chanY_n5  : std_ulogic := '0';
	signal track_4_1_chanY_n6  : std_ulogic := '0';
	signal track_4_1_chanY_n7  : std_ulogic := '0';
	signal track_4_1_chanY_n8  : std_ulogic := '0';
	signal track_4_1_chanY_n9  : std_ulogic := '0';
	signal track_4_2_chanX_n0  : std_ulogic := '0';
	signal track_4_2_chanX_n1  : std_ulogic := '0';
	signal track_4_2_chanX_n10 : std_ulogic := '0';
	signal track_4_2_chanX_n11 : std_ulogic := '0';
	signal track_4_2_chanX_n12 : std_ulogic := '0';
	signal track_4_2_chanX_n13 : std_ulogic := '0';
	signal track_4_2_chanX_n14 : std_ulogic := '0';
	signal track_4_2_chanX_n15 : std_ulogic := '0';
	signal track_4_2_chanX_n2  : std_ulogic := '0';
	signal track_4_2_chanX_n3  : std_ulogic := '0';
	signal track_4_2_chanX_n4  : std_ulogic := '0';
	signal track_4_2_chanX_n5  : std_ulogic := '0';
	signal track_4_2_chanX_n6  : std_ulogic := '0';
	signal track_4_2_chanX_n7  : std_ulogic := '0';
	signal track_4_2_chanX_n8  : std_ulogic := '0';
	signal track_4_2_chanX_n9  : std_ulogic := '0';
	signal track_4_2_chanY_n0  : std_ulogic := '0';
	signal track_4_2_chanY_n1  : std_ulogic := '0';
	signal track_4_2_chanY_n10 : std_ulogic := '0';
	signal track_4_2_chanY_n11 : std_ulogic := '0';
	signal track_4_2_chanY_n12 : std_ulogic := '0';
	signal track_4_2_chanY_n13 : std_ulogic := '0';
	signal track_4_2_chanY_n14 : std_ulogic := '0';
	signal track_4_2_chanY_n15 : std_ulogic := '0';
	signal track_4_2_chanY_n2  : std_ulogic := '0';
	signal track_4_2_chanY_n3  : std_ulogic := '0';
	signal track_4_2_chanY_n4  : std_ulogic := '0';
	signal track_4_2_chanY_n5  : std_ulogic := '0';
	signal track_4_2_chanY_n6  : std_ulogic := '0';
	signal track_4_2_chanY_n7  : std_ulogic := '0';
	signal track_4_2_chanY_n8  : std_ulogic := '0';
	signal track_4_2_chanY_n9  : std_ulogic := '0';
	signal track_4_3_chanX_n0  : std_ulogic := '0';
	signal track_4_3_chanX_n1  : std_ulogic := '0';
	signal track_4_3_chanX_n10 : std_ulogic := '0';
	signal track_4_3_chanX_n11 : std_ulogic := '0';
	signal track_4_3_chanX_n12 : std_ulogic := '0';
	signal track_4_3_chanX_n13 : std_ulogic := '0';
	signal track_4_3_chanX_n14 : std_ulogic := '0';
	signal track_4_3_chanX_n15 : std_ulogic := '0';
	signal track_4_3_chanX_n2  : std_ulogic := '0';
	signal track_4_3_chanX_n3  : std_ulogic := '0';
	signal track_4_3_chanX_n4  : std_ulogic := '0';
	signal track_4_3_chanX_n5  : std_ulogic := '0';
	signal track_4_3_chanX_n6  : std_ulogic := '0';
	signal track_4_3_chanX_n7  : std_ulogic := '0';
	signal track_4_3_chanX_n8  : std_ulogic := '0';
	signal track_4_3_chanX_n9  : std_ulogic := '0';
	signal track_4_3_chanY_n0  : std_ulogic := '0';
	signal track_4_3_chanY_n1  : std_ulogic := '0';
	signal track_4_3_chanY_n10 : std_ulogic := '0';
	signal track_4_3_chanY_n11 : std_ulogic := '0';
	signal track_4_3_chanY_n12 : std_ulogic := '0';
	signal track_4_3_chanY_n13 : std_ulogic := '0';
	signal track_4_3_chanY_n14 : std_ulogic := '0';
	signal track_4_3_chanY_n15 : std_ulogic := '0';
	signal track_4_3_chanY_n2  : std_ulogic := '0';
	signal track_4_3_chanY_n3  : std_ulogic := '0';
	signal track_4_3_chanY_n4  : std_ulogic := '0';
	signal track_4_3_chanY_n5  : std_ulogic := '0';
	signal track_4_3_chanY_n6  : std_ulogic := '0';
	signal track_4_3_chanY_n7  : std_ulogic := '0';
	signal track_4_3_chanY_n8  : std_ulogic := '0';
	signal track_4_3_chanY_n9  : std_ulogic := '0';
	signal track_4_4_chanX_n0  : std_ulogic := '0';
	signal track_4_4_chanX_n1  : std_ulogic := '0';
	signal track_4_4_chanX_n10 : std_ulogic := '0';
	signal track_4_4_chanX_n11 : std_ulogic := '0';
	signal track_4_4_chanX_n12 : std_ulogic := '0';
	signal track_4_4_chanX_n13 : std_ulogic := '0';
	signal track_4_4_chanX_n14 : std_ulogic := '0';
	signal track_4_4_chanX_n15 : std_ulogic := '0';
	signal track_4_4_chanX_n2  : std_ulogic := '0';
	signal track_4_4_chanX_n3  : std_ulogic := '0';
	signal track_4_4_chanX_n4  : std_ulogic := '0';
	signal track_4_4_chanX_n5  : std_ulogic := '0';
	signal track_4_4_chanX_n6  : std_ulogic := '0';
	signal track_4_4_chanX_n7  : std_ulogic := '0';
	signal track_4_4_chanX_n8  : std_ulogic := '0';
	signal track_4_4_chanX_n9  : std_ulogic := '0';
	signal track_4_4_chanY_n0  : std_ulogic := '0';
	signal track_4_4_chanY_n1  : std_ulogic := '0';
	signal track_4_4_chanY_n10 : std_ulogic := '0';
	signal track_4_4_chanY_n11 : std_ulogic := '0';
	signal track_4_4_chanY_n12 : std_ulogic := '0';
	signal track_4_4_chanY_n13 : std_ulogic := '0';
	signal track_4_4_chanY_n14 : std_ulogic := '0';
	signal track_4_4_chanY_n15 : std_ulogic := '0';
	signal track_4_4_chanY_n2  : std_ulogic := '0';
	signal track_4_4_chanY_n3  : std_ulogic := '0';
	signal track_4_4_chanY_n4  : std_ulogic := '0';
	signal track_4_4_chanY_n5  : std_ulogic := '0';
	signal track_4_4_chanY_n6  : std_ulogic := '0';
	signal track_4_4_chanY_n7  : std_ulogic := '0';
	signal track_4_4_chanY_n8  : std_ulogic := '0';
	signal track_4_4_chanY_n9  : std_ulogic := '0';
	signal track_4_5_chanX_n0  : std_ulogic := '0';
	signal track_4_5_chanX_n1  : std_ulogic := '0';
	signal track_4_5_chanX_n10 : std_ulogic := '0';
	signal track_4_5_chanX_n11 : std_ulogic := '0';
	signal track_4_5_chanX_n12 : std_ulogic := '0';
	signal track_4_5_chanX_n13 : std_ulogic := '0';
	signal track_4_5_chanX_n14 : std_ulogic := '0';
	signal track_4_5_chanX_n15 : std_ulogic := '0';
	signal track_4_5_chanX_n2  : std_ulogic := '0';
	signal track_4_5_chanX_n3  : std_ulogic := '0';
	signal track_4_5_chanX_n4  : std_ulogic := '0';
	signal track_4_5_chanX_n5  : std_ulogic := '0';
	signal track_4_5_chanX_n6  : std_ulogic := '0';
	signal track_4_5_chanX_n7  : std_ulogic := '0';
	signal track_4_5_chanX_n8  : std_ulogic := '0';
	signal track_4_5_chanX_n9  : std_ulogic := '0';
	signal track_4_5_chanY_n0  : std_ulogic := '0';
	signal track_4_5_chanY_n1  : std_ulogic := '0';
	signal track_4_5_chanY_n10 : std_ulogic := '0';
	signal track_4_5_chanY_n11 : std_ulogic := '0';
	signal track_4_5_chanY_n12 : std_ulogic := '0';
	signal track_4_5_chanY_n13 : std_ulogic := '0';
	signal track_4_5_chanY_n14 : std_ulogic := '0';
	signal track_4_5_chanY_n15 : std_ulogic := '0';
	signal track_4_5_chanY_n2  : std_ulogic := '0';
	signal track_4_5_chanY_n3  : std_ulogic := '0';
	signal track_4_5_chanY_n4  : std_ulogic := '0';
	signal track_4_5_chanY_n5  : std_ulogic := '0';
	signal track_4_5_chanY_n6  : std_ulogic := '0';
	signal track_4_5_chanY_n7  : std_ulogic := '0';
	signal track_4_5_chanY_n8  : std_ulogic := '0';
	signal track_4_5_chanY_n9  : std_ulogic := '0';
	signal track_4_6_chanX_n0  : std_ulogic := '0';
	signal track_4_6_chanX_n1  : std_ulogic := '0';
	signal track_4_6_chanX_n10 : std_ulogic := '0';
	signal track_4_6_chanX_n11 : std_ulogic := '0';
	signal track_4_6_chanX_n12 : std_ulogic := '0';
	signal track_4_6_chanX_n13 : std_ulogic := '0';
	signal track_4_6_chanX_n14 : std_ulogic := '0';
	signal track_4_6_chanX_n15 : std_ulogic := '0';
	signal track_4_6_chanX_n2  : std_ulogic := '0';
	signal track_4_6_chanX_n3  : std_ulogic := '0';
	signal track_4_6_chanX_n4  : std_ulogic := '0';
	signal track_4_6_chanX_n5  : std_ulogic := '0';
	signal track_4_6_chanX_n6  : std_ulogic := '0';
	signal track_4_6_chanX_n7  : std_ulogic := '0';
	signal track_4_6_chanX_n8  : std_ulogic := '0';
	signal track_4_6_chanX_n9  : std_ulogic := '0';
	signal track_4_6_chanY_n0  : std_ulogic := '0';
	signal track_4_6_chanY_n1  : std_ulogic := '0';
	signal track_4_6_chanY_n10 : std_ulogic := '0';
	signal track_4_6_chanY_n11 : std_ulogic := '0';
	signal track_4_6_chanY_n12 : std_ulogic := '0';
	signal track_4_6_chanY_n13 : std_ulogic := '0';
	signal track_4_6_chanY_n14 : std_ulogic := '0';
	signal track_4_6_chanY_n15 : std_ulogic := '0';
	signal track_4_6_chanY_n2  : std_ulogic := '0';
	signal track_4_6_chanY_n3  : std_ulogic := '0';
	signal track_4_6_chanY_n4  : std_ulogic := '0';
	signal track_4_6_chanY_n5  : std_ulogic := '0';
	signal track_4_6_chanY_n6  : std_ulogic := '0';
	signal track_4_6_chanY_n7  : std_ulogic := '0';
	signal track_4_6_chanY_n8  : std_ulogic := '0';
	signal track_4_6_chanY_n9  : std_ulogic := '0';
	signal track_5_0_chanX_n0  : std_ulogic := '0';
	signal track_5_0_chanX_n1  : std_ulogic := '0';
	signal track_5_0_chanX_n10 : std_ulogic := '0';
	signal track_5_0_chanX_n11 : std_ulogic := '0';
	signal track_5_0_chanX_n12 : std_ulogic := '0';
	signal track_5_0_chanX_n13 : std_ulogic := '0';
	signal track_5_0_chanX_n14 : std_ulogic := '0';
	signal track_5_0_chanX_n15 : std_ulogic := '0';
	signal track_5_0_chanX_n2  : std_ulogic := '0';
	signal track_5_0_chanX_n3  : std_ulogic := '0';
	signal track_5_0_chanX_n4  : std_ulogic := '0';
	signal track_5_0_chanX_n5  : std_ulogic := '0';
	signal track_5_0_chanX_n6  : std_ulogic := '0';
	signal track_5_0_chanX_n7  : std_ulogic := '0';
	signal track_5_0_chanX_n8  : std_ulogic := '0';
	signal track_5_0_chanX_n9  : std_ulogic := '0';
	signal track_5_1_chanX_n0  : std_ulogic := '0';
	signal track_5_1_chanX_n1  : std_ulogic := '0';
	signal track_5_1_chanX_n10 : std_ulogic := '0';
	signal track_5_1_chanX_n11 : std_ulogic := '0';
	signal track_5_1_chanX_n12 : std_ulogic := '0';
	signal track_5_1_chanX_n13 : std_ulogic := '0';
	signal track_5_1_chanX_n14 : std_ulogic := '0';
	signal track_5_1_chanX_n15 : std_ulogic := '0';
	signal track_5_1_chanX_n2  : std_ulogic := '0';
	signal track_5_1_chanX_n3  : std_ulogic := '0';
	signal track_5_1_chanX_n4  : std_ulogic := '0';
	signal track_5_1_chanX_n5  : std_ulogic := '0';
	signal track_5_1_chanX_n6  : std_ulogic := '0';
	signal track_5_1_chanX_n7  : std_ulogic := '0';
	signal track_5_1_chanX_n8  : std_ulogic := '0';
	signal track_5_1_chanX_n9  : std_ulogic := '0';
	signal track_5_1_chanY_n0  : std_ulogic := '0';
	signal track_5_1_chanY_n1  : std_ulogic := '0';
	signal track_5_1_chanY_n10 : std_ulogic := '0';
	signal track_5_1_chanY_n11 : std_ulogic := '0';
	signal track_5_1_chanY_n12 : std_ulogic := '0';
	signal track_5_1_chanY_n13 : std_ulogic := '0';
	signal track_5_1_chanY_n14 : std_ulogic := '0';
	signal track_5_1_chanY_n15 : std_ulogic := '0';
	signal track_5_1_chanY_n2  : std_ulogic := '0';
	signal track_5_1_chanY_n3  : std_ulogic := '0';
	signal track_5_1_chanY_n4  : std_ulogic := '0';
	signal track_5_1_chanY_n5  : std_ulogic := '0';
	signal track_5_1_chanY_n6  : std_ulogic := '0';
	signal track_5_1_chanY_n7  : std_ulogic := '0';
	signal track_5_1_chanY_n8  : std_ulogic := '0';
	signal track_5_1_chanY_n9  : std_ulogic := '0';
	signal track_5_2_chanX_n0  : std_ulogic := '0';
	signal track_5_2_chanX_n1  : std_ulogic := '0';
	signal track_5_2_chanX_n10 : std_ulogic := '0';
	signal track_5_2_chanX_n11 : std_ulogic := '0';
	signal track_5_2_chanX_n12 : std_ulogic := '0';
	signal track_5_2_chanX_n13 : std_ulogic := '0';
	signal track_5_2_chanX_n14 : std_ulogic := '0';
	signal track_5_2_chanX_n15 : std_ulogic := '0';
	signal track_5_2_chanX_n2  : std_ulogic := '0';
	signal track_5_2_chanX_n3  : std_ulogic := '0';
	signal track_5_2_chanX_n4  : std_ulogic := '0';
	signal track_5_2_chanX_n5  : std_ulogic := '0';
	signal track_5_2_chanX_n6  : std_ulogic := '0';
	signal track_5_2_chanX_n7  : std_ulogic := '0';
	signal track_5_2_chanX_n8  : std_ulogic := '0';
	signal track_5_2_chanX_n9  : std_ulogic := '0';
	signal track_5_2_chanY_n0  : std_ulogic := '0';
	signal track_5_2_chanY_n1  : std_ulogic := '0';
	signal track_5_2_chanY_n10 : std_ulogic := '0';
	signal track_5_2_chanY_n11 : std_ulogic := '0';
	signal track_5_2_chanY_n12 : std_ulogic := '0';
	signal track_5_2_chanY_n13 : std_ulogic := '0';
	signal track_5_2_chanY_n14 : std_ulogic := '0';
	signal track_5_2_chanY_n15 : std_ulogic := '0';
	signal track_5_2_chanY_n2  : std_ulogic := '0';
	signal track_5_2_chanY_n3  : std_ulogic := '0';
	signal track_5_2_chanY_n4  : std_ulogic := '0';
	signal track_5_2_chanY_n5  : std_ulogic := '0';
	signal track_5_2_chanY_n6  : std_ulogic := '0';
	signal track_5_2_chanY_n7  : std_ulogic := '0';
	signal track_5_2_chanY_n8  : std_ulogic := '0';
	signal track_5_2_chanY_n9  : std_ulogic := '0';
	signal track_5_3_chanX_n0  : std_ulogic := '0';
	signal track_5_3_chanX_n1  : std_ulogic := '0';
	signal track_5_3_chanX_n10 : std_ulogic := '0';
	signal track_5_3_chanX_n11 : std_ulogic := '0';
	signal track_5_3_chanX_n12 : std_ulogic := '0';
	signal track_5_3_chanX_n13 : std_ulogic := '0';
	signal track_5_3_chanX_n14 : std_ulogic := '0';
	signal track_5_3_chanX_n15 : std_ulogic := '0';
	signal track_5_3_chanX_n2  : std_ulogic := '0';
	signal track_5_3_chanX_n3  : std_ulogic := '0';
	signal track_5_3_chanX_n4  : std_ulogic := '0';
	signal track_5_3_chanX_n5  : std_ulogic := '0';
	signal track_5_3_chanX_n6  : std_ulogic := '0';
	signal track_5_3_chanX_n7  : std_ulogic := '0';
	signal track_5_3_chanX_n8  : std_ulogic := '0';
	signal track_5_3_chanX_n9  : std_ulogic := '0';
	signal track_5_3_chanY_n0  : std_ulogic := '0';
	signal track_5_3_chanY_n1  : std_ulogic := '0';
	signal track_5_3_chanY_n10 : std_ulogic := '0';
	signal track_5_3_chanY_n11 : std_ulogic := '0';
	signal track_5_3_chanY_n12 : std_ulogic := '0';
	signal track_5_3_chanY_n13 : std_ulogic := '0';
	signal track_5_3_chanY_n14 : std_ulogic := '0';
	signal track_5_3_chanY_n15 : std_ulogic := '0';
	signal track_5_3_chanY_n2  : std_ulogic := '0';
	signal track_5_3_chanY_n3  : std_ulogic := '0';
	signal track_5_3_chanY_n4  : std_ulogic := '0';
	signal track_5_3_chanY_n5  : std_ulogic := '0';
	signal track_5_3_chanY_n6  : std_ulogic := '0';
	signal track_5_3_chanY_n7  : std_ulogic := '0';
	signal track_5_3_chanY_n8  : std_ulogic := '0';
	signal track_5_3_chanY_n9  : std_ulogic := '0';
	signal track_5_4_chanX_n0  : std_ulogic := '0';
	signal track_5_4_chanX_n1  : std_ulogic := '0';
	signal track_5_4_chanX_n10 : std_ulogic := '0';
	signal track_5_4_chanX_n11 : std_ulogic := '0';
	signal track_5_4_chanX_n12 : std_ulogic := '0';
	signal track_5_4_chanX_n13 : std_ulogic := '0';
	signal track_5_4_chanX_n14 : std_ulogic := '0';
	signal track_5_4_chanX_n15 : std_ulogic := '0';
	signal track_5_4_chanX_n2  : std_ulogic := '0';
	signal track_5_4_chanX_n3  : std_ulogic := '0';
	signal track_5_4_chanX_n4  : std_ulogic := '0';
	signal track_5_4_chanX_n5  : std_ulogic := '0';
	signal track_5_4_chanX_n6  : std_ulogic := '0';
	signal track_5_4_chanX_n7  : std_ulogic := '0';
	signal track_5_4_chanX_n8  : std_ulogic := '0';
	signal track_5_4_chanX_n9  : std_ulogic := '0';
	signal track_5_4_chanY_n0  : std_ulogic := '0';
	signal track_5_4_chanY_n1  : std_ulogic := '0';
	signal track_5_4_chanY_n10 : std_ulogic := '0';
	signal track_5_4_chanY_n11 : std_ulogic := '0';
	signal track_5_4_chanY_n12 : std_ulogic := '0';
	signal track_5_4_chanY_n13 : std_ulogic := '0';
	signal track_5_4_chanY_n14 : std_ulogic := '0';
	signal track_5_4_chanY_n15 : std_ulogic := '0';
	signal track_5_4_chanY_n2  : std_ulogic := '0';
	signal track_5_4_chanY_n3  : std_ulogic := '0';
	signal track_5_4_chanY_n4  : std_ulogic := '0';
	signal track_5_4_chanY_n5  : std_ulogic := '0';
	signal track_5_4_chanY_n6  : std_ulogic := '0';
	signal track_5_4_chanY_n7  : std_ulogic := '0';
	signal track_5_4_chanY_n8  : std_ulogic := '0';
	signal track_5_4_chanY_n9  : std_ulogic := '0';
	signal track_5_5_chanX_n0  : std_ulogic := '0';
	signal track_5_5_chanX_n1  : std_ulogic := '0';
	signal track_5_5_chanX_n10 : std_ulogic := '0';
	signal track_5_5_chanX_n11 : std_ulogic := '0';
	signal track_5_5_chanX_n12 : std_ulogic := '0';
	signal track_5_5_chanX_n13 : std_ulogic := '0';
	signal track_5_5_chanX_n14 : std_ulogic := '0';
	signal track_5_5_chanX_n15 : std_ulogic := '0';
	signal track_5_5_chanX_n2  : std_ulogic := '0';
	signal track_5_5_chanX_n3  : std_ulogic := '0';
	signal track_5_5_chanX_n4  : std_ulogic := '0';
	signal track_5_5_chanX_n5  : std_ulogic := '0';
	signal track_5_5_chanX_n6  : std_ulogic := '0';
	signal track_5_5_chanX_n7  : std_ulogic := '0';
	signal track_5_5_chanX_n8  : std_ulogic := '0';
	signal track_5_5_chanX_n9  : std_ulogic := '0';
	signal track_5_5_chanY_n0  : std_ulogic := '0';
	signal track_5_5_chanY_n1  : std_ulogic := '0';
	signal track_5_5_chanY_n10 : std_ulogic := '0';
	signal track_5_5_chanY_n11 : std_ulogic := '0';
	signal track_5_5_chanY_n12 : std_ulogic := '0';
	signal track_5_5_chanY_n13 : std_ulogic := '0';
	signal track_5_5_chanY_n14 : std_ulogic := '0';
	signal track_5_5_chanY_n15 : std_ulogic := '0';
	signal track_5_5_chanY_n2  : std_ulogic := '0';
	signal track_5_5_chanY_n3  : std_ulogic := '0';
	signal track_5_5_chanY_n4  : std_ulogic := '0';
	signal track_5_5_chanY_n5  : std_ulogic := '0';
	signal track_5_5_chanY_n6  : std_ulogic := '0';
	signal track_5_5_chanY_n7  : std_ulogic := '0';
	signal track_5_5_chanY_n8  : std_ulogic := '0';
	signal track_5_5_chanY_n9  : std_ulogic := '0';
	signal track_5_6_chanX_n0  : std_ulogic := '0';
	signal track_5_6_chanX_n1  : std_ulogic := '0';
	signal track_5_6_chanX_n10 : std_ulogic := '0';
	signal track_5_6_chanX_n11 : std_ulogic := '0';
	signal track_5_6_chanX_n12 : std_ulogic := '0';
	signal track_5_6_chanX_n13 : std_ulogic := '0';
	signal track_5_6_chanX_n14 : std_ulogic := '0';
	signal track_5_6_chanX_n15 : std_ulogic := '0';
	signal track_5_6_chanX_n2  : std_ulogic := '0';
	signal track_5_6_chanX_n3  : std_ulogic := '0';
	signal track_5_6_chanX_n4  : std_ulogic := '0';
	signal track_5_6_chanX_n5  : std_ulogic := '0';
	signal track_5_6_chanX_n6  : std_ulogic := '0';
	signal track_5_6_chanX_n7  : std_ulogic := '0';
	signal track_5_6_chanX_n8  : std_ulogic := '0';
	signal track_5_6_chanX_n9  : std_ulogic := '0';
	signal track_5_6_chanY_n0  : std_ulogic := '0';
	signal track_5_6_chanY_n1  : std_ulogic := '0';
	signal track_5_6_chanY_n10 : std_ulogic := '0';
	signal track_5_6_chanY_n11 : std_ulogic := '0';
	signal track_5_6_chanY_n12 : std_ulogic := '0';
	signal track_5_6_chanY_n13 : std_ulogic := '0';
	signal track_5_6_chanY_n14 : std_ulogic := '0';
	signal track_5_6_chanY_n15 : std_ulogic := '0';
	signal track_5_6_chanY_n2  : std_ulogic := '0';
	signal track_5_6_chanY_n3  : std_ulogic := '0';
	signal track_5_6_chanY_n4  : std_ulogic := '0';
	signal track_5_6_chanY_n5  : std_ulogic := '0';
	signal track_5_6_chanY_n6  : std_ulogic := '0';
	signal track_5_6_chanY_n7  : std_ulogic := '0';
	signal track_5_6_chanY_n8  : std_ulogic := '0';
	signal track_5_6_chanY_n9  : std_ulogic := '0';
	signal track_6_0_chanX_n0  : std_ulogic := '0';
	signal track_6_0_chanX_n1  : std_ulogic := '0';
	signal track_6_0_chanX_n10 : std_ulogic := '0';
	signal track_6_0_chanX_n11 : std_ulogic := '0';
	signal track_6_0_chanX_n12 : std_ulogic := '0';
	signal track_6_0_chanX_n13 : std_ulogic := '0';
	signal track_6_0_chanX_n14 : std_ulogic := '0';
	signal track_6_0_chanX_n15 : std_ulogic := '0';
	signal track_6_0_chanX_n2  : std_ulogic := '0';
	signal track_6_0_chanX_n3  : std_ulogic := '0';
	signal track_6_0_chanX_n4  : std_ulogic := '0';
	signal track_6_0_chanX_n5  : std_ulogic := '0';
	signal track_6_0_chanX_n6  : std_ulogic := '0';
	signal track_6_0_chanX_n7  : std_ulogic := '0';
	signal track_6_0_chanX_n8  : std_ulogic := '0';
	signal track_6_0_chanX_n9  : std_ulogic := '0';
	signal track_6_1_chanX_n0  : std_ulogic := '0';
	signal track_6_1_chanX_n1  : std_ulogic := '0';
	signal track_6_1_chanX_n10 : std_ulogic := '0';
	signal track_6_1_chanX_n11 : std_ulogic := '0';
	signal track_6_1_chanX_n12 : std_ulogic := '0';
	signal track_6_1_chanX_n13 : std_ulogic := '0';
	signal track_6_1_chanX_n14 : std_ulogic := '0';
	signal track_6_1_chanX_n15 : std_ulogic := '0';
	signal track_6_1_chanX_n2  : std_ulogic := '0';
	signal track_6_1_chanX_n3  : std_ulogic := '0';
	signal track_6_1_chanX_n4  : std_ulogic := '0';
	signal track_6_1_chanX_n5  : std_ulogic := '0';
	signal track_6_1_chanX_n6  : std_ulogic := '0';
	signal track_6_1_chanX_n7  : std_ulogic := '0';
	signal track_6_1_chanX_n8  : std_ulogic := '0';
	signal track_6_1_chanX_n9  : std_ulogic := '0';
	signal track_6_1_chanY_n0  : std_ulogic := '0';
	signal track_6_1_chanY_n1  : std_ulogic := '0';
	signal track_6_1_chanY_n10 : std_ulogic := '0';
	signal track_6_1_chanY_n11 : std_ulogic := '0';
	signal track_6_1_chanY_n12 : std_ulogic := '0';
	signal track_6_1_chanY_n13 : std_ulogic := '0';
	signal track_6_1_chanY_n14 : std_ulogic := '0';
	signal track_6_1_chanY_n15 : std_ulogic := '0';
	signal track_6_1_chanY_n2  : std_ulogic := '0';
	signal track_6_1_chanY_n3  : std_ulogic := '0';
	signal track_6_1_chanY_n4  : std_ulogic := '0';
	signal track_6_1_chanY_n5  : std_ulogic := '0';
	signal track_6_1_chanY_n6  : std_ulogic := '0';
	signal track_6_1_chanY_n7  : std_ulogic := '0';
	signal track_6_1_chanY_n8  : std_ulogic := '0';
	signal track_6_1_chanY_n9  : std_ulogic := '0';
	signal track_6_2_chanX_n0  : std_ulogic := '0';
	signal track_6_2_chanX_n1  : std_ulogic := '0';
	signal track_6_2_chanX_n10 : std_ulogic := '0';
	signal track_6_2_chanX_n11 : std_ulogic := '0';
	signal track_6_2_chanX_n12 : std_ulogic := '0';
	signal track_6_2_chanX_n13 : std_ulogic := '0';
	signal track_6_2_chanX_n14 : std_ulogic := '0';
	signal track_6_2_chanX_n15 : std_ulogic := '0';
	signal track_6_2_chanX_n2  : std_ulogic := '0';
	signal track_6_2_chanX_n3  : std_ulogic := '0';
	signal track_6_2_chanX_n4  : std_ulogic := '0';
	signal track_6_2_chanX_n5  : std_ulogic := '0';
	signal track_6_2_chanX_n6  : std_ulogic := '0';
	signal track_6_2_chanX_n7  : std_ulogic := '0';
	signal track_6_2_chanX_n8  : std_ulogic := '0';
	signal track_6_2_chanX_n9  : std_ulogic := '0';
	signal track_6_2_chanY_n0  : std_ulogic := '0';
	signal track_6_2_chanY_n1  : std_ulogic := '0';
	signal track_6_2_chanY_n10 : std_ulogic := '0';
	signal track_6_2_chanY_n11 : std_ulogic := '0';
	signal track_6_2_chanY_n12 : std_ulogic := '0';
	signal track_6_2_chanY_n13 : std_ulogic := '0';
	signal track_6_2_chanY_n14 : std_ulogic := '0';
	signal track_6_2_chanY_n15 : std_ulogic := '0';
	signal track_6_2_chanY_n2  : std_ulogic := '0';
	signal track_6_2_chanY_n3  : std_ulogic := '0';
	signal track_6_2_chanY_n4  : std_ulogic := '0';
	signal track_6_2_chanY_n5  : std_ulogic := '0';
	signal track_6_2_chanY_n6  : std_ulogic := '0';
	signal track_6_2_chanY_n7  : std_ulogic := '0';
	signal track_6_2_chanY_n8  : std_ulogic := '0';
	signal track_6_2_chanY_n9  : std_ulogic := '0';
	signal track_6_3_chanX_n0  : std_ulogic := '0';
	signal track_6_3_chanX_n1  : std_ulogic := '0';
	signal track_6_3_chanX_n10 : std_ulogic := '0';
	signal track_6_3_chanX_n11 : std_ulogic := '0';
	signal track_6_3_chanX_n12 : std_ulogic := '0';
	signal track_6_3_chanX_n13 : std_ulogic := '0';
	signal track_6_3_chanX_n14 : std_ulogic := '0';
	signal track_6_3_chanX_n15 : std_ulogic := '0';
	signal track_6_3_chanX_n2  : std_ulogic := '0';
	signal track_6_3_chanX_n3  : std_ulogic := '0';
	signal track_6_3_chanX_n4  : std_ulogic := '0';
	signal track_6_3_chanX_n5  : std_ulogic := '0';
	signal track_6_3_chanX_n6  : std_ulogic := '0';
	signal track_6_3_chanX_n7  : std_ulogic := '0';
	signal track_6_3_chanX_n8  : std_ulogic := '0';
	signal track_6_3_chanX_n9  : std_ulogic := '0';
	signal track_6_3_chanY_n0  : std_ulogic := '0';
	signal track_6_3_chanY_n1  : std_ulogic := '0';
	signal track_6_3_chanY_n10 : std_ulogic := '0';
	signal track_6_3_chanY_n11 : std_ulogic := '0';
	signal track_6_3_chanY_n12 : std_ulogic := '0';
	signal track_6_3_chanY_n13 : std_ulogic := '0';
	signal track_6_3_chanY_n14 : std_ulogic := '0';
	signal track_6_3_chanY_n15 : std_ulogic := '0';
	signal track_6_3_chanY_n2  : std_ulogic := '0';
	signal track_6_3_chanY_n3  : std_ulogic := '0';
	signal track_6_3_chanY_n4  : std_ulogic := '0';
	signal track_6_3_chanY_n5  : std_ulogic := '0';
	signal track_6_3_chanY_n6  : std_ulogic := '0';
	signal track_6_3_chanY_n7  : std_ulogic := '0';
	signal track_6_3_chanY_n8  : std_ulogic := '0';
	signal track_6_3_chanY_n9  : std_ulogic := '0';
	signal track_6_4_chanX_n0  : std_ulogic := '0';
	signal track_6_4_chanX_n1  : std_ulogic := '0';
	signal track_6_4_chanX_n10 : std_ulogic := '0';
	signal track_6_4_chanX_n11 : std_ulogic := '0';
	signal track_6_4_chanX_n12 : std_ulogic := '0';
	signal track_6_4_chanX_n13 : std_ulogic := '0';
	signal track_6_4_chanX_n14 : std_ulogic := '0';
	signal track_6_4_chanX_n15 : std_ulogic := '0';
	signal track_6_4_chanX_n2  : std_ulogic := '0';
	signal track_6_4_chanX_n3  : std_ulogic := '0';
	signal track_6_4_chanX_n4  : std_ulogic := '0';
	signal track_6_4_chanX_n5  : std_ulogic := '0';
	signal track_6_4_chanX_n6  : std_ulogic := '0';
	signal track_6_4_chanX_n7  : std_ulogic := '0';
	signal track_6_4_chanX_n8  : std_ulogic := '0';
	signal track_6_4_chanX_n9  : std_ulogic := '0';
	signal track_6_4_chanY_n0  : std_ulogic := '0';
	signal track_6_4_chanY_n1  : std_ulogic := '0';
	signal track_6_4_chanY_n10 : std_ulogic := '0';
	signal track_6_4_chanY_n11 : std_ulogic := '0';
	signal track_6_4_chanY_n12 : std_ulogic := '0';
	signal track_6_4_chanY_n13 : std_ulogic := '0';
	signal track_6_4_chanY_n14 : std_ulogic := '0';
	signal track_6_4_chanY_n15 : std_ulogic := '0';
	signal track_6_4_chanY_n2  : std_ulogic := '0';
	signal track_6_4_chanY_n3  : std_ulogic := '0';
	signal track_6_4_chanY_n4  : std_ulogic := '0';
	signal track_6_4_chanY_n5  : std_ulogic := '0';
	signal track_6_4_chanY_n6  : std_ulogic := '0';
	signal track_6_4_chanY_n7  : std_ulogic := '0';
	signal track_6_4_chanY_n8  : std_ulogic := '0';
	signal track_6_4_chanY_n9  : std_ulogic := '0';
	signal track_6_5_chanX_n0  : std_ulogic := '0';
	signal track_6_5_chanX_n1  : std_ulogic := '0';
	signal track_6_5_chanX_n10 : std_ulogic := '0';
	signal track_6_5_chanX_n11 : std_ulogic := '0';
	signal track_6_5_chanX_n12 : std_ulogic := '0';
	signal track_6_5_chanX_n13 : std_ulogic := '0';
	signal track_6_5_chanX_n14 : std_ulogic := '0';
	signal track_6_5_chanX_n15 : std_ulogic := '0';
	signal track_6_5_chanX_n2  : std_ulogic := '0';
	signal track_6_5_chanX_n3  : std_ulogic := '0';
	signal track_6_5_chanX_n4  : std_ulogic := '0';
	signal track_6_5_chanX_n5  : std_ulogic := '0';
	signal track_6_5_chanX_n6  : std_ulogic := '0';
	signal track_6_5_chanX_n7  : std_ulogic := '0';
	signal track_6_5_chanX_n8  : std_ulogic := '0';
	signal track_6_5_chanX_n9  : std_ulogic := '0';
	signal track_6_5_chanY_n0  : std_ulogic := '0';
	signal track_6_5_chanY_n1  : std_ulogic := '0';
	signal track_6_5_chanY_n10 : std_ulogic := '0';
	signal track_6_5_chanY_n11 : std_ulogic := '0';
	signal track_6_5_chanY_n12 : std_ulogic := '0';
	signal track_6_5_chanY_n13 : std_ulogic := '0';
	signal track_6_5_chanY_n14 : std_ulogic := '0';
	signal track_6_5_chanY_n15 : std_ulogic := '0';
	signal track_6_5_chanY_n2  : std_ulogic := '0';
	signal track_6_5_chanY_n3  : std_ulogic := '0';
	signal track_6_5_chanY_n4  : std_ulogic := '0';
	signal track_6_5_chanY_n5  : std_ulogic := '0';
	signal track_6_5_chanY_n6  : std_ulogic := '0';
	signal track_6_5_chanY_n7  : std_ulogic := '0';
	signal track_6_5_chanY_n8  : std_ulogic := '0';
	signal track_6_5_chanY_n9  : std_ulogic := '0';
	signal track_6_6_chanX_n0  : std_ulogic := '0';
	signal track_6_6_chanX_n1  : std_ulogic := '0';
	signal track_6_6_chanX_n10 : std_ulogic := '0';
	signal track_6_6_chanX_n11 : std_ulogic := '0';
	signal track_6_6_chanX_n12 : std_ulogic := '0';
	signal track_6_6_chanX_n13 : std_ulogic := '0';
	signal track_6_6_chanX_n14 : std_ulogic := '0';
	signal track_6_6_chanX_n15 : std_ulogic := '0';
	signal track_6_6_chanX_n2  : std_ulogic := '0';
	signal track_6_6_chanX_n3  : std_ulogic := '0';
	signal track_6_6_chanX_n4  : std_ulogic := '0';
	signal track_6_6_chanX_n5  : std_ulogic := '0';
	signal track_6_6_chanX_n6  : std_ulogic := '0';
	signal track_6_6_chanX_n7  : std_ulogic := '0';
	signal track_6_6_chanX_n8  : std_ulogic := '0';
	signal track_6_6_chanX_n9  : std_ulogic := '0';
	signal track_6_6_chanY_n0  : std_ulogic := '0';
	signal track_6_6_chanY_n1  : std_ulogic := '0';
	signal track_6_6_chanY_n10 : std_ulogic := '0';
	signal track_6_6_chanY_n11 : std_ulogic := '0';
	signal track_6_6_chanY_n12 : std_ulogic := '0';
	signal track_6_6_chanY_n13 : std_ulogic := '0';
	signal track_6_6_chanY_n14 : std_ulogic := '0';
	signal track_6_6_chanY_n15 : std_ulogic := '0';
	signal track_6_6_chanY_n2  : std_ulogic := '0';
	signal track_6_6_chanY_n3  : std_ulogic := '0';
	signal track_6_6_chanY_n4  : std_ulogic := '0';
	signal track_6_6_chanY_n5  : std_ulogic := '0';
	signal track_6_6_chanY_n6  : std_ulogic := '0';
	signal track_6_6_chanY_n7  : std_ulogic := '0';
	signal track_6_6_chanY_n8  : std_ulogic := '0';
	signal track_6_6_chanY_n9  : std_ulogic := '0';
	signal track_7_0_chanX_n0  : std_ulogic := '0';
	signal track_7_0_chanX_n1  : std_ulogic := '0';
	signal track_7_0_chanX_n10 : std_ulogic := '0';
	signal track_7_0_chanX_n11 : std_ulogic := '0';
	signal track_7_0_chanX_n12 : std_ulogic := '0';
	signal track_7_0_chanX_n13 : std_ulogic := '0';
	signal track_7_0_chanX_n14 : std_ulogic := '0';
	signal track_7_0_chanX_n15 : std_ulogic := '0';
	signal track_7_0_chanX_n2  : std_ulogic := '0';
	signal track_7_0_chanX_n3  : std_ulogic := '0';
	signal track_7_0_chanX_n4  : std_ulogic := '0';
	signal track_7_0_chanX_n5  : std_ulogic := '0';
	signal track_7_0_chanX_n6  : std_ulogic := '0';
	signal track_7_0_chanX_n7  : std_ulogic := '0';
	signal track_7_0_chanX_n8  : std_ulogic := '0';
	signal track_7_0_chanX_n9  : std_ulogic := '0';
	signal track_7_1_chanX_n0  : std_ulogic := '0';
	signal track_7_1_chanX_n1  : std_ulogic := '0';
	signal track_7_1_chanX_n10 : std_ulogic := '0';
	signal track_7_1_chanX_n11 : std_ulogic := '0';
	signal track_7_1_chanX_n12 : std_ulogic := '0';
	signal track_7_1_chanX_n13 : std_ulogic := '0';
	signal track_7_1_chanX_n14 : std_ulogic := '0';
	signal track_7_1_chanX_n15 : std_ulogic := '0';
	signal track_7_1_chanX_n2  : std_ulogic := '0';
	signal track_7_1_chanX_n3  : std_ulogic := '0';
	signal track_7_1_chanX_n4  : std_ulogic := '0';
	signal track_7_1_chanX_n5  : std_ulogic := '0';
	signal track_7_1_chanX_n6  : std_ulogic := '0';
	signal track_7_1_chanX_n7  : std_ulogic := '0';
	signal track_7_1_chanX_n8  : std_ulogic := '0';
	signal track_7_1_chanX_n9  : std_ulogic := '0';
	signal track_7_1_chanY_n0  : std_ulogic := '0';
	signal track_7_1_chanY_n1  : std_ulogic := '0';
	signal track_7_1_chanY_n10 : std_ulogic := '0';
	signal track_7_1_chanY_n11 : std_ulogic := '0';
	signal track_7_1_chanY_n12 : std_ulogic := '0';
	signal track_7_1_chanY_n13 : std_ulogic := '0';
	signal track_7_1_chanY_n14 : std_ulogic := '0';
	signal track_7_1_chanY_n15 : std_ulogic := '0';
	signal track_7_1_chanY_n2  : std_ulogic := '0';
	signal track_7_1_chanY_n3  : std_ulogic := '0';
	signal track_7_1_chanY_n4  : std_ulogic := '0';
	signal track_7_1_chanY_n5  : std_ulogic := '0';
	signal track_7_1_chanY_n6  : std_ulogic := '0';
	signal track_7_1_chanY_n7  : std_ulogic := '0';
	signal track_7_1_chanY_n8  : std_ulogic := '0';
	signal track_7_1_chanY_n9  : std_ulogic := '0';
	signal track_7_2_chanX_n0  : std_ulogic := '0';
	signal track_7_2_chanX_n1  : std_ulogic := '0';
	signal track_7_2_chanX_n10 : std_ulogic := '0';
	signal track_7_2_chanX_n11 : std_ulogic := '0';
	signal track_7_2_chanX_n12 : std_ulogic := '0';
	signal track_7_2_chanX_n13 : std_ulogic := '0';
	signal track_7_2_chanX_n14 : std_ulogic := '0';
	signal track_7_2_chanX_n15 : std_ulogic := '0';
	signal track_7_2_chanX_n2  : std_ulogic := '0';
	signal track_7_2_chanX_n3  : std_ulogic := '0';
	signal track_7_2_chanX_n4  : std_ulogic := '0';
	signal track_7_2_chanX_n5  : std_ulogic := '0';
	signal track_7_2_chanX_n6  : std_ulogic := '0';
	signal track_7_2_chanX_n7  : std_ulogic := '0';
	signal track_7_2_chanX_n8  : std_ulogic := '0';
	signal track_7_2_chanX_n9  : std_ulogic := '0';
	signal track_7_2_chanY_n0  : std_ulogic := '0';
	signal track_7_2_chanY_n1  : std_ulogic := '0';
	signal track_7_2_chanY_n10 : std_ulogic := '0';
	signal track_7_2_chanY_n11 : std_ulogic := '0';
	signal track_7_2_chanY_n12 : std_ulogic := '0';
	signal track_7_2_chanY_n13 : std_ulogic := '0';
	signal track_7_2_chanY_n14 : std_ulogic := '0';
	signal track_7_2_chanY_n15 : std_ulogic := '0';
	signal track_7_2_chanY_n2  : std_ulogic := '0';
	signal track_7_2_chanY_n3  : std_ulogic := '0';
	signal track_7_2_chanY_n4  : std_ulogic := '0';
	signal track_7_2_chanY_n5  : std_ulogic := '0';
	signal track_7_2_chanY_n6  : std_ulogic := '0';
	signal track_7_2_chanY_n7  : std_ulogic := '0';
	signal track_7_2_chanY_n8  : std_ulogic := '0';
	signal track_7_2_chanY_n9  : std_ulogic := '0';
	signal track_7_3_chanX_n0  : std_ulogic := '0';
	signal track_7_3_chanX_n1  : std_ulogic := '0';
	signal track_7_3_chanX_n10 : std_ulogic := '0';
	signal track_7_3_chanX_n11 : std_ulogic := '0';
	signal track_7_3_chanX_n12 : std_ulogic := '0';
	signal track_7_3_chanX_n13 : std_ulogic := '0';
	signal track_7_3_chanX_n14 : std_ulogic := '0';
	signal track_7_3_chanX_n15 : std_ulogic := '0';
	signal track_7_3_chanX_n2  : std_ulogic := '0';
	signal track_7_3_chanX_n3  : std_ulogic := '0';
	signal track_7_3_chanX_n4  : std_ulogic := '0';
	signal track_7_3_chanX_n5  : std_ulogic := '0';
	signal track_7_3_chanX_n6  : std_ulogic := '0';
	signal track_7_3_chanX_n7  : std_ulogic := '0';
	signal track_7_3_chanX_n8  : std_ulogic := '0';
	signal track_7_3_chanX_n9  : std_ulogic := '0';
	signal track_7_3_chanY_n0  : std_ulogic := '0';
	signal track_7_3_chanY_n1  : std_ulogic := '0';
	signal track_7_3_chanY_n10 : std_ulogic := '0';
	signal track_7_3_chanY_n11 : std_ulogic := '0';
	signal track_7_3_chanY_n12 : std_ulogic := '0';
	signal track_7_3_chanY_n13 : std_ulogic := '0';
	signal track_7_3_chanY_n14 : std_ulogic := '0';
	signal track_7_3_chanY_n15 : std_ulogic := '0';
	signal track_7_3_chanY_n2  : std_ulogic := '0';
	signal track_7_3_chanY_n3  : std_ulogic := '0';
	signal track_7_3_chanY_n4  : std_ulogic := '0';
	signal track_7_3_chanY_n5  : std_ulogic := '0';
	signal track_7_3_chanY_n6  : std_ulogic := '0';
	signal track_7_3_chanY_n7  : std_ulogic := '0';
	signal track_7_3_chanY_n8  : std_ulogic := '0';
	signal track_7_3_chanY_n9  : std_ulogic := '0';
	signal track_7_4_chanX_n0  : std_ulogic := '0';
	signal track_7_4_chanX_n1  : std_ulogic := '0';
	signal track_7_4_chanX_n10 : std_ulogic := '0';
	signal track_7_4_chanX_n11 : std_ulogic := '0';
	signal track_7_4_chanX_n12 : std_ulogic := '0';
	signal track_7_4_chanX_n13 : std_ulogic := '0';
	signal track_7_4_chanX_n14 : std_ulogic := '0';
	signal track_7_4_chanX_n15 : std_ulogic := '0';
	signal track_7_4_chanX_n2  : std_ulogic := '0';
	signal track_7_4_chanX_n3  : std_ulogic := '0';
	signal track_7_4_chanX_n4  : std_ulogic := '0';
	signal track_7_4_chanX_n5  : std_ulogic := '0';
	signal track_7_4_chanX_n6  : std_ulogic := '0';
	signal track_7_4_chanX_n7  : std_ulogic := '0';
	signal track_7_4_chanX_n8  : std_ulogic := '0';
	signal track_7_4_chanX_n9  : std_ulogic := '0';
	signal track_7_4_chanY_n0  : std_ulogic := '0';
	signal track_7_4_chanY_n1  : std_ulogic := '0';
	signal track_7_4_chanY_n10 : std_ulogic := '0';
	signal track_7_4_chanY_n11 : std_ulogic := '0';
	signal track_7_4_chanY_n12 : std_ulogic := '0';
	signal track_7_4_chanY_n13 : std_ulogic := '0';
	signal track_7_4_chanY_n14 : std_ulogic := '0';
	signal track_7_4_chanY_n15 : std_ulogic := '0';
	signal track_7_4_chanY_n2  : std_ulogic := '0';
	signal track_7_4_chanY_n3  : std_ulogic := '0';
	signal track_7_4_chanY_n4  : std_ulogic := '0';
	signal track_7_4_chanY_n5  : std_ulogic := '0';
	signal track_7_4_chanY_n6  : std_ulogic := '0';
	signal track_7_4_chanY_n7  : std_ulogic := '0';
	signal track_7_4_chanY_n8  : std_ulogic := '0';
	signal track_7_4_chanY_n9  : std_ulogic := '0';
	signal track_7_5_chanX_n0  : std_ulogic := '0';
	signal track_7_5_chanX_n1  : std_ulogic := '0';
	signal track_7_5_chanX_n10 : std_ulogic := '0';
	signal track_7_5_chanX_n11 : std_ulogic := '0';
	signal track_7_5_chanX_n12 : std_ulogic := '0';
	signal track_7_5_chanX_n13 : std_ulogic := '0';
	signal track_7_5_chanX_n14 : std_ulogic := '0';
	signal track_7_5_chanX_n15 : std_ulogic := '0';
	signal track_7_5_chanX_n2  : std_ulogic := '0';
	signal track_7_5_chanX_n3  : std_ulogic := '0';
	signal track_7_5_chanX_n4  : std_ulogic := '0';
	signal track_7_5_chanX_n5  : std_ulogic := '0';
	signal track_7_5_chanX_n6  : std_ulogic := '0';
	signal track_7_5_chanX_n7  : std_ulogic := '0';
	signal track_7_5_chanX_n8  : std_ulogic := '0';
	signal track_7_5_chanX_n9  : std_ulogic := '0';
	signal track_7_5_chanY_n0  : std_ulogic := '0';
	signal track_7_5_chanY_n1  : std_ulogic := '0';
	signal track_7_5_chanY_n10 : std_ulogic := '0';
	signal track_7_5_chanY_n11 : std_ulogic := '0';
	signal track_7_5_chanY_n12 : std_ulogic := '0';
	signal track_7_5_chanY_n13 : std_ulogic := '0';
	signal track_7_5_chanY_n14 : std_ulogic := '0';
	signal track_7_5_chanY_n15 : std_ulogic := '0';
	signal track_7_5_chanY_n2  : std_ulogic := '0';
	signal track_7_5_chanY_n3  : std_ulogic := '0';
	signal track_7_5_chanY_n4  : std_ulogic := '0';
	signal track_7_5_chanY_n5  : std_ulogic := '0';
	signal track_7_5_chanY_n6  : std_ulogic := '0';
	signal track_7_5_chanY_n7  : std_ulogic := '0';
	signal track_7_5_chanY_n8  : std_ulogic := '0';
	signal track_7_5_chanY_n9  : std_ulogic := '0';
	signal track_7_6_chanX_n0  : std_ulogic := '0';
	signal track_7_6_chanX_n1  : std_ulogic := '0';
	signal track_7_6_chanX_n10 : std_ulogic := '0';
	signal track_7_6_chanX_n11 : std_ulogic := '0';
	signal track_7_6_chanX_n12 : std_ulogic := '0';
	signal track_7_6_chanX_n13 : std_ulogic := '0';
	signal track_7_6_chanX_n14 : std_ulogic := '0';
	signal track_7_6_chanX_n15 : std_ulogic := '0';
	signal track_7_6_chanX_n2  : std_ulogic := '0';
	signal track_7_6_chanX_n3  : std_ulogic := '0';
	signal track_7_6_chanX_n4  : std_ulogic := '0';
	signal track_7_6_chanX_n5  : std_ulogic := '0';
	signal track_7_6_chanX_n6  : std_ulogic := '0';
	signal track_7_6_chanX_n7  : std_ulogic := '0';
	signal track_7_6_chanX_n8  : std_ulogic := '0';
	signal track_7_6_chanX_n9  : std_ulogic := '0';
	signal track_7_6_chanY_n0  : std_ulogic := '0';
	signal track_7_6_chanY_n1  : std_ulogic := '0';
	signal track_7_6_chanY_n10 : std_ulogic := '0';
	signal track_7_6_chanY_n11 : std_ulogic := '0';
	signal track_7_6_chanY_n12 : std_ulogic := '0';
	signal track_7_6_chanY_n13 : std_ulogic := '0';
	signal track_7_6_chanY_n14 : std_ulogic := '0';
	signal track_7_6_chanY_n15 : std_ulogic := '0';
	signal track_7_6_chanY_n2  : std_ulogic := '0';
	signal track_7_6_chanY_n3  : std_ulogic := '0';
	signal track_7_6_chanY_n4  : std_ulogic := '0';
	signal track_7_6_chanY_n5  : std_ulogic := '0';
	signal track_7_6_chanY_n6  : std_ulogic := '0';
	signal track_7_6_chanY_n7  : std_ulogic := '0';
	signal track_7_6_chanY_n8  : std_ulogic := '0';
	signal track_7_6_chanY_n9  : std_ulogic := '0';
	signal track_8_0_chanX_n0  : std_ulogic := '0';
	signal track_8_0_chanX_n1  : std_ulogic := '0';
	signal track_8_0_chanX_n10 : std_ulogic := '0';
	signal track_8_0_chanX_n11 : std_ulogic := '0';
	signal track_8_0_chanX_n12 : std_ulogic := '0';
	signal track_8_0_chanX_n13 : std_ulogic := '0';
	signal track_8_0_chanX_n14 : std_ulogic := '0';
	signal track_8_0_chanX_n15 : std_ulogic := '0';
	signal track_8_0_chanX_n2  : std_ulogic := '0';
	signal track_8_0_chanX_n3  : std_ulogic := '0';
	signal track_8_0_chanX_n4  : std_ulogic := '0';
	signal track_8_0_chanX_n5  : std_ulogic := '0';
	signal track_8_0_chanX_n6  : std_ulogic := '0';
	signal track_8_0_chanX_n7  : std_ulogic := '0';
	signal track_8_0_chanX_n8  : std_ulogic := '0';
	signal track_8_0_chanX_n9  : std_ulogic := '0';
	signal track_8_1_chanX_n0  : std_ulogic := '0';
	signal track_8_1_chanX_n1  : std_ulogic := '0';
	signal track_8_1_chanX_n10 : std_ulogic := '0';
	signal track_8_1_chanX_n11 : std_ulogic := '0';
	signal track_8_1_chanX_n12 : std_ulogic := '0';
	signal track_8_1_chanX_n13 : std_ulogic := '0';
	signal track_8_1_chanX_n14 : std_ulogic := '0';
	signal track_8_1_chanX_n15 : std_ulogic := '0';
	signal track_8_1_chanX_n2  : std_ulogic := '0';
	signal track_8_1_chanX_n3  : std_ulogic := '0';
	signal track_8_1_chanX_n4  : std_ulogic := '0';
	signal track_8_1_chanX_n5  : std_ulogic := '0';
	signal track_8_1_chanX_n6  : std_ulogic := '0';
	signal track_8_1_chanX_n7  : std_ulogic := '0';
	signal track_8_1_chanX_n8  : std_ulogic := '0';
	signal track_8_1_chanX_n9  : std_ulogic := '0';
	signal track_8_1_chanY_n0  : std_ulogic := '0';
	signal track_8_1_chanY_n1  : std_ulogic := '0';
	signal track_8_1_chanY_n10 : std_ulogic := '0';
	signal track_8_1_chanY_n11 : std_ulogic := '0';
	signal track_8_1_chanY_n12 : std_ulogic := '0';
	signal track_8_1_chanY_n13 : std_ulogic := '0';
	signal track_8_1_chanY_n14 : std_ulogic := '0';
	signal track_8_1_chanY_n15 : std_ulogic := '0';
	signal track_8_1_chanY_n2  : std_ulogic := '0';
	signal track_8_1_chanY_n3  : std_ulogic := '0';
	signal track_8_1_chanY_n4  : std_ulogic := '0';
	signal track_8_1_chanY_n5  : std_ulogic := '0';
	signal track_8_1_chanY_n6  : std_ulogic := '0';
	signal track_8_1_chanY_n7  : std_ulogic := '0';
	signal track_8_1_chanY_n8  : std_ulogic := '0';
	signal track_8_1_chanY_n9  : std_ulogic := '0';
	signal track_8_2_chanX_n0  : std_ulogic := '0';
	signal track_8_2_chanX_n1  : std_ulogic := '0';
	signal track_8_2_chanX_n10 : std_ulogic := '0';
	signal track_8_2_chanX_n11 : std_ulogic := '0';
	signal track_8_2_chanX_n12 : std_ulogic := '0';
	signal track_8_2_chanX_n13 : std_ulogic := '0';
	signal track_8_2_chanX_n14 : std_ulogic := '0';
	signal track_8_2_chanX_n15 : std_ulogic := '0';
	signal track_8_2_chanX_n2  : std_ulogic := '0';
	signal track_8_2_chanX_n3  : std_ulogic := '0';
	signal track_8_2_chanX_n4  : std_ulogic := '0';
	signal track_8_2_chanX_n5  : std_ulogic := '0';
	signal track_8_2_chanX_n6  : std_ulogic := '0';
	signal track_8_2_chanX_n7  : std_ulogic := '0';
	signal track_8_2_chanX_n8  : std_ulogic := '0';
	signal track_8_2_chanX_n9  : std_ulogic := '0';
	signal track_8_2_chanY_n0  : std_ulogic := '0';
	signal track_8_2_chanY_n1  : std_ulogic := '0';
	signal track_8_2_chanY_n10 : std_ulogic := '0';
	signal track_8_2_chanY_n11 : std_ulogic := '0';
	signal track_8_2_chanY_n12 : std_ulogic := '0';
	signal track_8_2_chanY_n13 : std_ulogic := '0';
	signal track_8_2_chanY_n14 : std_ulogic := '0';
	signal track_8_2_chanY_n15 : std_ulogic := '0';
	signal track_8_2_chanY_n2  : std_ulogic := '0';
	signal track_8_2_chanY_n3  : std_ulogic := '0';
	signal track_8_2_chanY_n4  : std_ulogic := '0';
	signal track_8_2_chanY_n5  : std_ulogic := '0';
	signal track_8_2_chanY_n6  : std_ulogic := '0';
	signal track_8_2_chanY_n7  : std_ulogic := '0';
	signal track_8_2_chanY_n8  : std_ulogic := '0';
	signal track_8_2_chanY_n9  : std_ulogic := '0';
	signal track_8_3_chanX_n0  : std_ulogic := '0';
	signal track_8_3_chanX_n1  : std_ulogic := '0';
	signal track_8_3_chanX_n10 : std_ulogic := '0';
	signal track_8_3_chanX_n11 : std_ulogic := '0';
	signal track_8_3_chanX_n12 : std_ulogic := '0';
	signal track_8_3_chanX_n13 : std_ulogic := '0';
	signal track_8_3_chanX_n14 : std_ulogic := '0';
	signal track_8_3_chanX_n15 : std_ulogic := '0';
	signal track_8_3_chanX_n2  : std_ulogic := '0';
	signal track_8_3_chanX_n3  : std_ulogic := '0';
	signal track_8_3_chanX_n4  : std_ulogic := '0';
	signal track_8_3_chanX_n5  : std_ulogic := '0';
	signal track_8_3_chanX_n6  : std_ulogic := '0';
	signal track_8_3_chanX_n7  : std_ulogic := '0';
	signal track_8_3_chanX_n8  : std_ulogic := '0';
	signal track_8_3_chanX_n9  : std_ulogic := '0';
	signal track_8_3_chanY_n0  : std_ulogic := '0';
	signal track_8_3_chanY_n1  : std_ulogic := '0';
	signal track_8_3_chanY_n10 : std_ulogic := '0';
	signal track_8_3_chanY_n11 : std_ulogic := '0';
	signal track_8_3_chanY_n12 : std_ulogic := '0';
	signal track_8_3_chanY_n13 : std_ulogic := '0';
	signal track_8_3_chanY_n14 : std_ulogic := '0';
	signal track_8_3_chanY_n15 : std_ulogic := '0';
	signal track_8_3_chanY_n2  : std_ulogic := '0';
	signal track_8_3_chanY_n3  : std_ulogic := '0';
	signal track_8_3_chanY_n4  : std_ulogic := '0';
	signal track_8_3_chanY_n5  : std_ulogic := '0';
	signal track_8_3_chanY_n6  : std_ulogic := '0';
	signal track_8_3_chanY_n7  : std_ulogic := '0';
	signal track_8_3_chanY_n8  : std_ulogic := '0';
	signal track_8_3_chanY_n9  : std_ulogic := '0';
	signal track_8_4_chanX_n0  : std_ulogic := '0';
	signal track_8_4_chanX_n1  : std_ulogic := '0';
	signal track_8_4_chanX_n10 : std_ulogic := '0';
	signal track_8_4_chanX_n11 : std_ulogic := '0';
	signal track_8_4_chanX_n12 : std_ulogic := '0';
	signal track_8_4_chanX_n13 : std_ulogic := '0';
	signal track_8_4_chanX_n14 : std_ulogic := '0';
	signal track_8_4_chanX_n15 : std_ulogic := '0';
	signal track_8_4_chanX_n2  : std_ulogic := '0';
	signal track_8_4_chanX_n3  : std_ulogic := '0';
	signal track_8_4_chanX_n4  : std_ulogic := '0';
	signal track_8_4_chanX_n5  : std_ulogic := '0';
	signal track_8_4_chanX_n6  : std_ulogic := '0';
	signal track_8_4_chanX_n7  : std_ulogic := '0';
	signal track_8_4_chanX_n8  : std_ulogic := '0';
	signal track_8_4_chanX_n9  : std_ulogic := '0';
	signal track_8_4_chanY_n0  : std_ulogic := '0';
	signal track_8_4_chanY_n1  : std_ulogic := '0';
	signal track_8_4_chanY_n10 : std_ulogic := '0';
	signal track_8_4_chanY_n11 : std_ulogic := '0';
	signal track_8_4_chanY_n12 : std_ulogic := '0';
	signal track_8_4_chanY_n13 : std_ulogic := '0';
	signal track_8_4_chanY_n14 : std_ulogic := '0';
	signal track_8_4_chanY_n15 : std_ulogic := '0';
	signal track_8_4_chanY_n2  : std_ulogic := '0';
	signal track_8_4_chanY_n3  : std_ulogic := '0';
	signal track_8_4_chanY_n4  : std_ulogic := '0';
	signal track_8_4_chanY_n5  : std_ulogic := '0';
	signal track_8_4_chanY_n6  : std_ulogic := '0';
	signal track_8_4_chanY_n7  : std_ulogic := '0';
	signal track_8_4_chanY_n8  : std_ulogic := '0';
	signal track_8_4_chanY_n9  : std_ulogic := '0';
	signal track_8_5_chanX_n0  : std_ulogic := '0';
	signal track_8_5_chanX_n1  : std_ulogic := '0';
	signal track_8_5_chanX_n10 : std_ulogic := '0';
	signal track_8_5_chanX_n11 : std_ulogic := '0';
	signal track_8_5_chanX_n12 : std_ulogic := '0';
	signal track_8_5_chanX_n13 : std_ulogic := '0';
	signal track_8_5_chanX_n14 : std_ulogic := '0';
	signal track_8_5_chanX_n15 : std_ulogic := '0';
	signal track_8_5_chanX_n2  : std_ulogic := '0';
	signal track_8_5_chanX_n3  : std_ulogic := '0';
	signal track_8_5_chanX_n4  : std_ulogic := '0';
	signal track_8_5_chanX_n5  : std_ulogic := '0';
	signal track_8_5_chanX_n6  : std_ulogic := '0';
	signal track_8_5_chanX_n7  : std_ulogic := '0';
	signal track_8_5_chanX_n8  : std_ulogic := '0';
	signal track_8_5_chanX_n9  : std_ulogic := '0';
	signal track_8_5_chanY_n0  : std_ulogic := '0';
	signal track_8_5_chanY_n1  : std_ulogic := '0';
	signal track_8_5_chanY_n10 : std_ulogic := '0';
	signal track_8_5_chanY_n11 : std_ulogic := '0';
	signal track_8_5_chanY_n12 : std_ulogic := '0';
	signal track_8_5_chanY_n13 : std_ulogic := '0';
	signal track_8_5_chanY_n14 : std_ulogic := '0';
	signal track_8_5_chanY_n15 : std_ulogic := '0';
	signal track_8_5_chanY_n2  : std_ulogic := '0';
	signal track_8_5_chanY_n3  : std_ulogic := '0';
	signal track_8_5_chanY_n4  : std_ulogic := '0';
	signal track_8_5_chanY_n5  : std_ulogic := '0';
	signal track_8_5_chanY_n6  : std_ulogic := '0';
	signal track_8_5_chanY_n7  : std_ulogic := '0';
	signal track_8_5_chanY_n8  : std_ulogic := '0';
	signal track_8_5_chanY_n9  : std_ulogic := '0';
	signal track_8_6_chanX_n0  : std_ulogic := '0';
	signal track_8_6_chanX_n1  : std_ulogic := '0';
	signal track_8_6_chanX_n10 : std_ulogic := '0';
	signal track_8_6_chanX_n11 : std_ulogic := '0';
	signal track_8_6_chanX_n12 : std_ulogic := '0';
	signal track_8_6_chanX_n13 : std_ulogic := '0';
	signal track_8_6_chanX_n14 : std_ulogic := '0';
	signal track_8_6_chanX_n15 : std_ulogic := '0';
	signal track_8_6_chanX_n2  : std_ulogic := '0';
	signal track_8_6_chanX_n3  : std_ulogic := '0';
	signal track_8_6_chanX_n4  : std_ulogic := '0';
	signal track_8_6_chanX_n5  : std_ulogic := '0';
	signal track_8_6_chanX_n6  : std_ulogic := '0';
	signal track_8_6_chanX_n7  : std_ulogic := '0';
	signal track_8_6_chanX_n8  : std_ulogic := '0';
	signal track_8_6_chanX_n9  : std_ulogic := '0';
	signal track_8_6_chanY_n0  : std_ulogic := '0';
	signal track_8_6_chanY_n1  : std_ulogic := '0';
	signal track_8_6_chanY_n10 : std_ulogic := '0';
	signal track_8_6_chanY_n11 : std_ulogic := '0';
	signal track_8_6_chanY_n12 : std_ulogic := '0';
	signal track_8_6_chanY_n13 : std_ulogic := '0';
	signal track_8_6_chanY_n14 : std_ulogic := '0';
	signal track_8_6_chanY_n15 : std_ulogic := '0';
	signal track_8_6_chanY_n2  : std_ulogic := '0';
	signal track_8_6_chanY_n3  : std_ulogic := '0';
	signal track_8_6_chanY_n4  : std_ulogic := '0';
	signal track_8_6_chanY_n5  : std_ulogic := '0';
	signal track_8_6_chanY_n6  : std_ulogic := '0';
	signal track_8_6_chanY_n7  : std_ulogic := '0';
	signal track_8_6_chanY_n8  : std_ulogic := '0';
	signal track_8_6_chanY_n9  : std_ulogic := '0';

	-- Input pins fanin choices (inputs of the mux driving the pin) --
	signal CLB_1_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_0_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_1_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_2_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_3_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_4_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_5_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_6_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_7_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_8_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_IN_pin_9_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal IO_0_1_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_1_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_2_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_2_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_3_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_3_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_4_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_4_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_5_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_5_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_6_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_0_6_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_1_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_1_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_1_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_1_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_2_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_2_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_2_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_2_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_3_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_3_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_3_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_3_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_4_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_4_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_4_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_4_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_5_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_5_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_5_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_5_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_6_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_6_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_6_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_6_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_7_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_7_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_7_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_7_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_8_0_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_8_0_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_8_7_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_8_7_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_1_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_1_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_2_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_2_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_3_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_3_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_4_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_4_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_5_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_5_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_6_IN_pin_0_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');
	signal IO_9_6_IN_pin_1_driver_mux_fanins  : std_ulogic_vector(7 downto 0) := (others => '0');

	-- Input pins selectors (selector of the mux driving the pin, i.e. the bitstream portion configuring the input pin) --
	signal CLB_1_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_1_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_2_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_3_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_4_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_5_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_6_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_7_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_1_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_2_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_3_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_4_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_5_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_0_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_1_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_2_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_3_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_4_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_5_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_6_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_7_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_8_driver_mux_selector : integer range 0 to 3 := 0;
	signal CLB_8_6_IN_pin_9_driver_mux_selector : integer range 0 to 3 := 0;
	signal IO_0_1_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_1_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_2_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_2_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_3_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_3_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_4_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_4_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_5_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_5_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_6_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_0_6_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_1_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_1_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_1_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_1_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_2_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_2_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_2_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_2_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_3_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_3_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_3_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_3_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_4_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_4_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_4_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_4_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_5_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_5_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_5_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_5_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_6_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_6_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_6_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_6_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_7_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_7_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_7_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_7_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_8_0_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_8_0_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_8_7_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_8_7_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_1_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_1_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_2_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_2_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_3_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_3_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_4_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_4_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_5_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_5_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_6_IN_pin_0_driver_mux_selector  : integer range 0 to 7 := 0;
	signal IO_9_6_IN_pin_1_driver_mux_selector  : integer range 0 to 7 := 0;

	-- Tracks fanin choices (inputs of the mux driving the track) --
	signal track_0_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_0_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_0_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_1_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_1_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_2_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_3_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_4_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_5_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_6_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_7_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n11_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_0_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n13_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_0_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n15_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_0_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_0_chanX_n9_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_1_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n10_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_1_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n12_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_1_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n14_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_1_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_1_chanY_n8_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_1_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_2_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_3_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_4_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanX_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n11_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n13_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n15_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_5_chanY_n9_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n11_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanX_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n13_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanX_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n15_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanX_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanX_n9_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanY_n0_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n1_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n10_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n11_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanY_n12_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n13_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanY_n14_driver_mux_fanins : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n15_driver_mux_fanins : std_ulogic_vector(1 downto 0) := (others => '0');
	signal track_8_6_chanY_n2_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n3_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n4_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n5_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n6_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n7_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n8_driver_mux_fanins  : std_ulogic_vector(3 downto 0) := (others => '0');
	signal track_8_6_chanY_n9_driver_mux_fanins  : std_ulogic_vector(1 downto 0) := (others => '0');

	-- Tracks selectors (selector of the mux driving the track, i.e. the bitstream portion configuring the track) --
	signal track_0_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n10_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n12_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n14_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_1_chanY_n8_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_0_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n11_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n13_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n15_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_0_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_0_6_chanY_n9_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_1_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n10_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n12_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n14_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_0_chanX_n8_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_1_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n10_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n12_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n14_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_1_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanX_n8_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_1_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_1_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_2_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_3_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_4_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_5_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_6_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_0_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_7_6_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n11_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_0_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n13_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_0_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n15_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_0_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_0_chanX_n9_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_8_1_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n10_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_1_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n12_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_1_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n14_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_1_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_1_chanY_n8_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_8_1_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_2_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_3_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_4_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanX_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n11_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n13_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n15_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_5_chanY_n9_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n11_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanX_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n13_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanX_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n15_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanX_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanX_n9_driver_mux_selector  : integer range 0 to 1 := 0;
	signal track_8_6_chanY_n0_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n1_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n10_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n11_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanY_n12_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n13_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanY_n14_driver_mux_selector : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n15_driver_mux_selector : integer range 0 to 1 := 0;
	signal track_8_6_chanY_n2_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n3_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n4_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n5_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n6_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n7_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n8_driver_mux_selector  : integer range 0 to 3 := 0;
	signal track_8_6_chanY_n9_driver_mux_selector  : integer range 0 to 1 := 0;

	-- CLB inputs --
	signal CLB_1_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_1_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_1_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_1_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_1_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_1_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_2_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_3_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_4_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_5_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_6_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_7_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_1_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_2_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_3_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_4_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_5_inputs : std_ulogic_vector(9 downto 0) := (others => '0');
	signal CLB_8_6_inputs : std_ulogic_vector(9 downto 0) := (others => '0');

	-- CLB outputs --
	signal CLB_1_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_outputs : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_outputs : std_ulogic_vector(3 downto 0) := (others => '0');

	-- CLB snapshot out --
	signal CLB_1_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_1_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_2_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_3_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_4_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_5_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_6_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_7_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_1_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_2_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_3_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_4_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_5_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');
	signal CLB_8_6_snapshot_out : std_ulogic_vector(3 downto 0) := (others => '0');

begin

	-- Input pins fanin choices (inputs of the mux driving the pin) --
	CLB_1_1_IN_pin_0_driver_mux_fanins <= track_1_1_chanX_n9 & track_1_1_chanX_n8 & track_1_1_chanX_n1 & track_1_1_chanX_n0;
	CLB_1_1_IN_pin_1_driver_mux_fanins <= track_1_1_chanY_n9 & track_1_1_chanY_n8 & track_1_1_chanY_n1 & track_1_1_chanY_n0;
	CLB_1_1_IN_pin_2_driver_mux_fanins <= track_1_0_chanX_n9 & track_1_0_chanX_n8 & track_1_0_chanX_n1 & track_1_0_chanX_n0;
	CLB_1_1_IN_pin_3_driver_mux_fanins <= track_0_1_chanY_n11 & track_0_1_chanY_n10 & track_0_1_chanY_n3 & track_0_1_chanY_n2;
	CLB_1_1_IN_pin_4_driver_mux_fanins <= track_1_1_chanX_n11 & track_1_1_chanX_n10 & track_1_1_chanX_n3 & track_1_1_chanX_n2;
	CLB_1_1_IN_pin_5_driver_mux_fanins <= track_1_1_chanY_n13 & track_1_1_chanY_n12 & track_1_1_chanY_n5 & track_1_1_chanY_n4;
	CLB_1_1_IN_pin_6_driver_mux_fanins <= track_1_0_chanX_n13 & track_1_0_chanX_n12 & track_1_0_chanX_n5 & track_1_0_chanX_n4;
	CLB_1_1_IN_pin_7_driver_mux_fanins <= track_0_1_chanY_n13 & track_0_1_chanY_n12 & track_0_1_chanY_n5 & track_0_1_chanY_n4;
	CLB_1_1_IN_pin_8_driver_mux_fanins <= track_1_1_chanX_n15 & track_1_1_chanX_n14 & track_1_1_chanX_n7 & track_1_1_chanX_n6;
	CLB_1_1_IN_pin_9_driver_mux_fanins <= track_1_1_chanY_n15 & track_1_1_chanY_n14 & track_1_1_chanY_n7 & track_1_1_chanY_n6;
	CLB_1_2_IN_pin_0_driver_mux_fanins <= track_1_2_chanX_n9 & track_1_2_chanX_n8 & track_1_2_chanX_n1 & track_1_2_chanX_n0;
	CLB_1_2_IN_pin_1_driver_mux_fanins <= track_1_2_chanY_n9 & track_1_2_chanY_n8 & track_1_2_chanY_n1 & track_1_2_chanY_n0;
	CLB_1_2_IN_pin_2_driver_mux_fanins <= track_1_1_chanX_n9 & track_1_1_chanX_n8 & track_1_1_chanX_n1 & track_1_1_chanX_n0;
	CLB_1_2_IN_pin_3_driver_mux_fanins <= track_0_2_chanY_n11 & track_0_2_chanY_n10 & track_0_2_chanY_n3 & track_0_2_chanY_n2;
	CLB_1_2_IN_pin_4_driver_mux_fanins <= track_1_2_chanX_n11 & track_1_2_chanX_n10 & track_1_2_chanX_n3 & track_1_2_chanX_n2;
	CLB_1_2_IN_pin_5_driver_mux_fanins <= track_1_2_chanY_n13 & track_1_2_chanY_n12 & track_1_2_chanY_n5 & track_1_2_chanY_n4;
	CLB_1_2_IN_pin_6_driver_mux_fanins <= track_1_1_chanX_n13 & track_1_1_chanX_n12 & track_1_1_chanX_n5 & track_1_1_chanX_n4;
	CLB_1_2_IN_pin_7_driver_mux_fanins <= track_0_2_chanY_n13 & track_0_2_chanY_n12 & track_0_2_chanY_n5 & track_0_2_chanY_n4;
	CLB_1_2_IN_pin_8_driver_mux_fanins <= track_1_2_chanX_n15 & track_1_2_chanX_n14 & track_1_2_chanX_n7 & track_1_2_chanX_n6;
	CLB_1_2_IN_pin_9_driver_mux_fanins <= track_1_2_chanY_n15 & track_1_2_chanY_n14 & track_1_2_chanY_n7 & track_1_2_chanY_n6;
	CLB_1_3_IN_pin_0_driver_mux_fanins <= track_1_3_chanX_n9 & track_1_3_chanX_n8 & track_1_3_chanX_n1 & track_1_3_chanX_n0;
	CLB_1_3_IN_pin_1_driver_mux_fanins <= track_1_3_chanY_n9 & track_1_3_chanY_n8 & track_1_3_chanY_n1 & track_1_3_chanY_n0;
	CLB_1_3_IN_pin_2_driver_mux_fanins <= track_1_2_chanX_n9 & track_1_2_chanX_n8 & track_1_2_chanX_n1 & track_1_2_chanX_n0;
	CLB_1_3_IN_pin_3_driver_mux_fanins <= track_0_3_chanY_n11 & track_0_3_chanY_n10 & track_0_3_chanY_n3 & track_0_3_chanY_n2;
	CLB_1_3_IN_pin_4_driver_mux_fanins <= track_1_3_chanX_n11 & track_1_3_chanX_n10 & track_1_3_chanX_n3 & track_1_3_chanX_n2;
	CLB_1_3_IN_pin_5_driver_mux_fanins <= track_1_3_chanY_n13 & track_1_3_chanY_n12 & track_1_3_chanY_n5 & track_1_3_chanY_n4;
	CLB_1_3_IN_pin_6_driver_mux_fanins <= track_1_2_chanX_n13 & track_1_2_chanX_n12 & track_1_2_chanX_n5 & track_1_2_chanX_n4;
	CLB_1_3_IN_pin_7_driver_mux_fanins <= track_0_3_chanY_n13 & track_0_3_chanY_n12 & track_0_3_chanY_n5 & track_0_3_chanY_n4;
	CLB_1_3_IN_pin_8_driver_mux_fanins <= track_1_3_chanX_n15 & track_1_3_chanX_n14 & track_1_3_chanX_n7 & track_1_3_chanX_n6;
	CLB_1_3_IN_pin_9_driver_mux_fanins <= track_1_3_chanY_n15 & track_1_3_chanY_n14 & track_1_3_chanY_n7 & track_1_3_chanY_n6;
	CLB_1_4_IN_pin_0_driver_mux_fanins <= track_1_4_chanX_n9 & track_1_4_chanX_n8 & track_1_4_chanX_n1 & track_1_4_chanX_n0;
	CLB_1_4_IN_pin_1_driver_mux_fanins <= track_1_4_chanY_n9 & track_1_4_chanY_n8 & track_1_4_chanY_n1 & track_1_4_chanY_n0;
	CLB_1_4_IN_pin_2_driver_mux_fanins <= track_1_3_chanX_n9 & track_1_3_chanX_n8 & track_1_3_chanX_n1 & track_1_3_chanX_n0;
	CLB_1_4_IN_pin_3_driver_mux_fanins <= track_0_4_chanY_n11 & track_0_4_chanY_n10 & track_0_4_chanY_n3 & track_0_4_chanY_n2;
	CLB_1_4_IN_pin_4_driver_mux_fanins <= track_1_4_chanX_n11 & track_1_4_chanX_n10 & track_1_4_chanX_n3 & track_1_4_chanX_n2;
	CLB_1_4_IN_pin_5_driver_mux_fanins <= track_1_4_chanY_n13 & track_1_4_chanY_n12 & track_1_4_chanY_n5 & track_1_4_chanY_n4;
	CLB_1_4_IN_pin_6_driver_mux_fanins <= track_1_3_chanX_n13 & track_1_3_chanX_n12 & track_1_3_chanX_n5 & track_1_3_chanX_n4;
	CLB_1_4_IN_pin_7_driver_mux_fanins <= track_0_4_chanY_n13 & track_0_4_chanY_n12 & track_0_4_chanY_n5 & track_0_4_chanY_n4;
	CLB_1_4_IN_pin_8_driver_mux_fanins <= track_1_4_chanX_n15 & track_1_4_chanX_n14 & track_1_4_chanX_n7 & track_1_4_chanX_n6;
	CLB_1_4_IN_pin_9_driver_mux_fanins <= track_1_4_chanY_n15 & track_1_4_chanY_n14 & track_1_4_chanY_n7 & track_1_4_chanY_n6;
	CLB_1_5_IN_pin_0_driver_mux_fanins <= track_1_5_chanX_n9 & track_1_5_chanX_n8 & track_1_5_chanX_n1 & track_1_5_chanX_n0;
	CLB_1_5_IN_pin_1_driver_mux_fanins <= track_1_5_chanY_n9 & track_1_5_chanY_n8 & track_1_5_chanY_n1 & track_1_5_chanY_n0;
	CLB_1_5_IN_pin_2_driver_mux_fanins <= track_1_4_chanX_n9 & track_1_4_chanX_n8 & track_1_4_chanX_n1 & track_1_4_chanX_n0;
	CLB_1_5_IN_pin_3_driver_mux_fanins <= track_0_5_chanY_n11 & track_0_5_chanY_n10 & track_0_5_chanY_n3 & track_0_5_chanY_n2;
	CLB_1_5_IN_pin_4_driver_mux_fanins <= track_1_5_chanX_n11 & track_1_5_chanX_n10 & track_1_5_chanX_n3 & track_1_5_chanX_n2;
	CLB_1_5_IN_pin_5_driver_mux_fanins <= track_1_5_chanY_n13 & track_1_5_chanY_n12 & track_1_5_chanY_n5 & track_1_5_chanY_n4;
	CLB_1_5_IN_pin_6_driver_mux_fanins <= track_1_4_chanX_n13 & track_1_4_chanX_n12 & track_1_4_chanX_n5 & track_1_4_chanX_n4;
	CLB_1_5_IN_pin_7_driver_mux_fanins <= track_0_5_chanY_n13 & track_0_5_chanY_n12 & track_0_5_chanY_n5 & track_0_5_chanY_n4;
	CLB_1_5_IN_pin_8_driver_mux_fanins <= track_1_5_chanX_n15 & track_1_5_chanX_n14 & track_1_5_chanX_n7 & track_1_5_chanX_n6;
	CLB_1_5_IN_pin_9_driver_mux_fanins <= track_1_5_chanY_n15 & track_1_5_chanY_n14 & track_1_5_chanY_n7 & track_1_5_chanY_n6;
	CLB_1_6_IN_pin_0_driver_mux_fanins <= track_1_6_chanX_n9 & track_1_6_chanX_n8 & track_1_6_chanX_n1 & track_1_6_chanX_n0;
	CLB_1_6_IN_pin_1_driver_mux_fanins <= track_1_6_chanY_n9 & track_1_6_chanY_n8 & track_1_6_chanY_n1 & track_1_6_chanY_n0;
	CLB_1_6_IN_pin_2_driver_mux_fanins <= track_1_5_chanX_n9 & track_1_5_chanX_n8 & track_1_5_chanX_n1 & track_1_5_chanX_n0;
	CLB_1_6_IN_pin_3_driver_mux_fanins <= track_0_6_chanY_n11 & track_0_6_chanY_n10 & track_0_6_chanY_n3 & track_0_6_chanY_n2;
	CLB_1_6_IN_pin_4_driver_mux_fanins <= track_1_6_chanX_n11 & track_1_6_chanX_n10 & track_1_6_chanX_n3 & track_1_6_chanX_n2;
	CLB_1_6_IN_pin_5_driver_mux_fanins <= track_1_6_chanY_n13 & track_1_6_chanY_n12 & track_1_6_chanY_n5 & track_1_6_chanY_n4;
	CLB_1_6_IN_pin_6_driver_mux_fanins <= track_1_5_chanX_n13 & track_1_5_chanX_n12 & track_1_5_chanX_n5 & track_1_5_chanX_n4;
	CLB_1_6_IN_pin_7_driver_mux_fanins <= track_0_6_chanY_n13 & track_0_6_chanY_n12 & track_0_6_chanY_n5 & track_0_6_chanY_n4;
	CLB_1_6_IN_pin_8_driver_mux_fanins <= track_1_6_chanX_n15 & track_1_6_chanX_n14 & track_1_6_chanX_n7 & track_1_6_chanX_n6;
	CLB_1_6_IN_pin_9_driver_mux_fanins <= track_1_6_chanY_n15 & track_1_6_chanY_n14 & track_1_6_chanY_n7 & track_1_6_chanY_n6;
	CLB_2_1_IN_pin_0_driver_mux_fanins <= track_2_1_chanX_n9 & track_2_1_chanX_n8 & track_2_1_chanX_n1 & track_2_1_chanX_n0;
	CLB_2_1_IN_pin_1_driver_mux_fanins <= track_2_1_chanY_n9 & track_2_1_chanY_n8 & track_2_1_chanY_n1 & track_2_1_chanY_n0;
	CLB_2_1_IN_pin_2_driver_mux_fanins <= track_2_0_chanX_n9 & track_2_0_chanX_n8 & track_2_0_chanX_n1 & track_2_0_chanX_n0;
	CLB_2_1_IN_pin_3_driver_mux_fanins <= track_1_1_chanY_n11 & track_1_1_chanY_n10 & track_1_1_chanY_n3 & track_1_1_chanY_n2;
	CLB_2_1_IN_pin_4_driver_mux_fanins <= track_2_1_chanX_n11 & track_2_1_chanX_n10 & track_2_1_chanX_n3 & track_2_1_chanX_n2;
	CLB_2_1_IN_pin_5_driver_mux_fanins <= track_2_1_chanY_n13 & track_2_1_chanY_n12 & track_2_1_chanY_n5 & track_2_1_chanY_n4;
	CLB_2_1_IN_pin_6_driver_mux_fanins <= track_2_0_chanX_n13 & track_2_0_chanX_n12 & track_2_0_chanX_n5 & track_2_0_chanX_n4;
	CLB_2_1_IN_pin_7_driver_mux_fanins <= track_1_1_chanY_n13 & track_1_1_chanY_n12 & track_1_1_chanY_n5 & track_1_1_chanY_n4;
	CLB_2_1_IN_pin_8_driver_mux_fanins <= track_2_1_chanX_n15 & track_2_1_chanX_n14 & track_2_1_chanX_n7 & track_2_1_chanX_n6;
	CLB_2_1_IN_pin_9_driver_mux_fanins <= track_2_1_chanY_n15 & track_2_1_chanY_n14 & track_2_1_chanY_n7 & track_2_1_chanY_n6;
	CLB_2_2_IN_pin_0_driver_mux_fanins <= track_2_2_chanX_n9 & track_2_2_chanX_n8 & track_2_2_chanX_n1 & track_2_2_chanX_n0;
	CLB_2_2_IN_pin_1_driver_mux_fanins <= track_2_2_chanY_n9 & track_2_2_chanY_n8 & track_2_2_chanY_n1 & track_2_2_chanY_n0;
	CLB_2_2_IN_pin_2_driver_mux_fanins <= track_2_1_chanX_n9 & track_2_1_chanX_n8 & track_2_1_chanX_n1 & track_2_1_chanX_n0;
	CLB_2_2_IN_pin_3_driver_mux_fanins <= track_1_2_chanY_n11 & track_1_2_chanY_n10 & track_1_2_chanY_n3 & track_1_2_chanY_n2;
	CLB_2_2_IN_pin_4_driver_mux_fanins <= track_2_2_chanX_n11 & track_2_2_chanX_n10 & track_2_2_chanX_n3 & track_2_2_chanX_n2;
	CLB_2_2_IN_pin_5_driver_mux_fanins <= track_2_2_chanY_n13 & track_2_2_chanY_n12 & track_2_2_chanY_n5 & track_2_2_chanY_n4;
	CLB_2_2_IN_pin_6_driver_mux_fanins <= track_2_1_chanX_n13 & track_2_1_chanX_n12 & track_2_1_chanX_n5 & track_2_1_chanX_n4;
	CLB_2_2_IN_pin_7_driver_mux_fanins <= track_1_2_chanY_n13 & track_1_2_chanY_n12 & track_1_2_chanY_n5 & track_1_2_chanY_n4;
	CLB_2_2_IN_pin_8_driver_mux_fanins <= track_2_2_chanX_n15 & track_2_2_chanX_n14 & track_2_2_chanX_n7 & track_2_2_chanX_n6;
	CLB_2_2_IN_pin_9_driver_mux_fanins <= track_2_2_chanY_n15 & track_2_2_chanY_n14 & track_2_2_chanY_n7 & track_2_2_chanY_n6;
	CLB_2_3_IN_pin_0_driver_mux_fanins <= track_2_3_chanX_n9 & track_2_3_chanX_n8 & track_2_3_chanX_n1 & track_2_3_chanX_n0;
	CLB_2_3_IN_pin_1_driver_mux_fanins <= track_2_3_chanY_n9 & track_2_3_chanY_n8 & track_2_3_chanY_n1 & track_2_3_chanY_n0;
	CLB_2_3_IN_pin_2_driver_mux_fanins <= track_2_2_chanX_n9 & track_2_2_chanX_n8 & track_2_2_chanX_n1 & track_2_2_chanX_n0;
	CLB_2_3_IN_pin_3_driver_mux_fanins <= track_1_3_chanY_n11 & track_1_3_chanY_n10 & track_1_3_chanY_n3 & track_1_3_chanY_n2;
	CLB_2_3_IN_pin_4_driver_mux_fanins <= track_2_3_chanX_n11 & track_2_3_chanX_n10 & track_2_3_chanX_n3 & track_2_3_chanX_n2;
	CLB_2_3_IN_pin_5_driver_mux_fanins <= track_2_3_chanY_n13 & track_2_3_chanY_n12 & track_2_3_chanY_n5 & track_2_3_chanY_n4;
	CLB_2_3_IN_pin_6_driver_mux_fanins <= track_2_2_chanX_n13 & track_2_2_chanX_n12 & track_2_2_chanX_n5 & track_2_2_chanX_n4;
	CLB_2_3_IN_pin_7_driver_mux_fanins <= track_1_3_chanY_n13 & track_1_3_chanY_n12 & track_1_3_chanY_n5 & track_1_3_chanY_n4;
	CLB_2_3_IN_pin_8_driver_mux_fanins <= track_2_3_chanX_n15 & track_2_3_chanX_n14 & track_2_3_chanX_n7 & track_2_3_chanX_n6;
	CLB_2_3_IN_pin_9_driver_mux_fanins <= track_2_3_chanY_n15 & track_2_3_chanY_n14 & track_2_3_chanY_n7 & track_2_3_chanY_n6;
	CLB_2_4_IN_pin_0_driver_mux_fanins <= track_2_4_chanX_n9 & track_2_4_chanX_n8 & track_2_4_chanX_n1 & track_2_4_chanX_n0;
	CLB_2_4_IN_pin_1_driver_mux_fanins <= track_2_4_chanY_n9 & track_2_4_chanY_n8 & track_2_4_chanY_n1 & track_2_4_chanY_n0;
	CLB_2_4_IN_pin_2_driver_mux_fanins <= track_2_3_chanX_n9 & track_2_3_chanX_n8 & track_2_3_chanX_n1 & track_2_3_chanX_n0;
	CLB_2_4_IN_pin_3_driver_mux_fanins <= track_1_4_chanY_n11 & track_1_4_chanY_n10 & track_1_4_chanY_n3 & track_1_4_chanY_n2;
	CLB_2_4_IN_pin_4_driver_mux_fanins <= track_2_4_chanX_n11 & track_2_4_chanX_n10 & track_2_4_chanX_n3 & track_2_4_chanX_n2;
	CLB_2_4_IN_pin_5_driver_mux_fanins <= track_2_4_chanY_n13 & track_2_4_chanY_n12 & track_2_4_chanY_n5 & track_2_4_chanY_n4;
	CLB_2_4_IN_pin_6_driver_mux_fanins <= track_2_3_chanX_n13 & track_2_3_chanX_n12 & track_2_3_chanX_n5 & track_2_3_chanX_n4;
	CLB_2_4_IN_pin_7_driver_mux_fanins <= track_1_4_chanY_n13 & track_1_4_chanY_n12 & track_1_4_chanY_n5 & track_1_4_chanY_n4;
	CLB_2_4_IN_pin_8_driver_mux_fanins <= track_2_4_chanX_n15 & track_2_4_chanX_n14 & track_2_4_chanX_n7 & track_2_4_chanX_n6;
	CLB_2_4_IN_pin_9_driver_mux_fanins <= track_2_4_chanY_n15 & track_2_4_chanY_n14 & track_2_4_chanY_n7 & track_2_4_chanY_n6;
	CLB_2_5_IN_pin_0_driver_mux_fanins <= track_2_5_chanX_n9 & track_2_5_chanX_n8 & track_2_5_chanX_n1 & track_2_5_chanX_n0;
	CLB_2_5_IN_pin_1_driver_mux_fanins <= track_2_5_chanY_n9 & track_2_5_chanY_n8 & track_2_5_chanY_n1 & track_2_5_chanY_n0;
	CLB_2_5_IN_pin_2_driver_mux_fanins <= track_2_4_chanX_n9 & track_2_4_chanX_n8 & track_2_4_chanX_n1 & track_2_4_chanX_n0;
	CLB_2_5_IN_pin_3_driver_mux_fanins <= track_1_5_chanY_n11 & track_1_5_chanY_n10 & track_1_5_chanY_n3 & track_1_5_chanY_n2;
	CLB_2_5_IN_pin_4_driver_mux_fanins <= track_2_5_chanX_n11 & track_2_5_chanX_n10 & track_2_5_chanX_n3 & track_2_5_chanX_n2;
	CLB_2_5_IN_pin_5_driver_mux_fanins <= track_2_5_chanY_n13 & track_2_5_chanY_n12 & track_2_5_chanY_n5 & track_2_5_chanY_n4;
	CLB_2_5_IN_pin_6_driver_mux_fanins <= track_2_4_chanX_n13 & track_2_4_chanX_n12 & track_2_4_chanX_n5 & track_2_4_chanX_n4;
	CLB_2_5_IN_pin_7_driver_mux_fanins <= track_1_5_chanY_n13 & track_1_5_chanY_n12 & track_1_5_chanY_n5 & track_1_5_chanY_n4;
	CLB_2_5_IN_pin_8_driver_mux_fanins <= track_2_5_chanX_n15 & track_2_5_chanX_n14 & track_2_5_chanX_n7 & track_2_5_chanX_n6;
	CLB_2_5_IN_pin_9_driver_mux_fanins <= track_2_5_chanY_n15 & track_2_5_chanY_n14 & track_2_5_chanY_n7 & track_2_5_chanY_n6;
	CLB_2_6_IN_pin_0_driver_mux_fanins <= track_2_6_chanX_n9 & track_2_6_chanX_n8 & track_2_6_chanX_n1 & track_2_6_chanX_n0;
	CLB_2_6_IN_pin_1_driver_mux_fanins <= track_2_6_chanY_n9 & track_2_6_chanY_n8 & track_2_6_chanY_n1 & track_2_6_chanY_n0;
	CLB_2_6_IN_pin_2_driver_mux_fanins <= track_2_5_chanX_n9 & track_2_5_chanX_n8 & track_2_5_chanX_n1 & track_2_5_chanX_n0;
	CLB_2_6_IN_pin_3_driver_mux_fanins <= track_1_6_chanY_n11 & track_1_6_chanY_n10 & track_1_6_chanY_n3 & track_1_6_chanY_n2;
	CLB_2_6_IN_pin_4_driver_mux_fanins <= track_2_6_chanX_n11 & track_2_6_chanX_n10 & track_2_6_chanX_n3 & track_2_6_chanX_n2;
	CLB_2_6_IN_pin_5_driver_mux_fanins <= track_2_6_chanY_n13 & track_2_6_chanY_n12 & track_2_6_chanY_n5 & track_2_6_chanY_n4;
	CLB_2_6_IN_pin_6_driver_mux_fanins <= track_2_5_chanX_n13 & track_2_5_chanX_n12 & track_2_5_chanX_n5 & track_2_5_chanX_n4;
	CLB_2_6_IN_pin_7_driver_mux_fanins <= track_1_6_chanY_n13 & track_1_6_chanY_n12 & track_1_6_chanY_n5 & track_1_6_chanY_n4;
	CLB_2_6_IN_pin_8_driver_mux_fanins <= track_2_6_chanX_n15 & track_2_6_chanX_n14 & track_2_6_chanX_n7 & track_2_6_chanX_n6;
	CLB_2_6_IN_pin_9_driver_mux_fanins <= track_2_6_chanY_n15 & track_2_6_chanY_n14 & track_2_6_chanY_n7 & track_2_6_chanY_n6;
	CLB_3_1_IN_pin_0_driver_mux_fanins <= track_3_1_chanX_n9 & track_3_1_chanX_n8 & track_3_1_chanX_n1 & track_3_1_chanX_n0;
	CLB_3_1_IN_pin_1_driver_mux_fanins <= track_3_1_chanY_n9 & track_3_1_chanY_n8 & track_3_1_chanY_n1 & track_3_1_chanY_n0;
	CLB_3_1_IN_pin_2_driver_mux_fanins <= track_3_0_chanX_n9 & track_3_0_chanX_n8 & track_3_0_chanX_n1 & track_3_0_chanX_n0;
	CLB_3_1_IN_pin_3_driver_mux_fanins <= track_2_1_chanY_n11 & track_2_1_chanY_n10 & track_2_1_chanY_n3 & track_2_1_chanY_n2;
	CLB_3_1_IN_pin_4_driver_mux_fanins <= track_3_1_chanX_n11 & track_3_1_chanX_n10 & track_3_1_chanX_n3 & track_3_1_chanX_n2;
	CLB_3_1_IN_pin_5_driver_mux_fanins <= track_3_1_chanY_n13 & track_3_1_chanY_n12 & track_3_1_chanY_n5 & track_3_1_chanY_n4;
	CLB_3_1_IN_pin_6_driver_mux_fanins <= track_3_0_chanX_n13 & track_3_0_chanX_n12 & track_3_0_chanX_n5 & track_3_0_chanX_n4;
	CLB_3_1_IN_pin_7_driver_mux_fanins <= track_2_1_chanY_n13 & track_2_1_chanY_n12 & track_2_1_chanY_n5 & track_2_1_chanY_n4;
	CLB_3_1_IN_pin_8_driver_mux_fanins <= track_3_1_chanX_n15 & track_3_1_chanX_n14 & track_3_1_chanX_n7 & track_3_1_chanX_n6;
	CLB_3_1_IN_pin_9_driver_mux_fanins <= track_3_1_chanY_n15 & track_3_1_chanY_n14 & track_3_1_chanY_n7 & track_3_1_chanY_n6;
	CLB_3_2_IN_pin_0_driver_mux_fanins <= track_3_2_chanX_n9 & track_3_2_chanX_n8 & track_3_2_chanX_n1 & track_3_2_chanX_n0;
	CLB_3_2_IN_pin_1_driver_mux_fanins <= track_3_2_chanY_n9 & track_3_2_chanY_n8 & track_3_2_chanY_n1 & track_3_2_chanY_n0;
	CLB_3_2_IN_pin_2_driver_mux_fanins <= track_3_1_chanX_n9 & track_3_1_chanX_n8 & track_3_1_chanX_n1 & track_3_1_chanX_n0;
	CLB_3_2_IN_pin_3_driver_mux_fanins <= track_2_2_chanY_n11 & track_2_2_chanY_n10 & track_2_2_chanY_n3 & track_2_2_chanY_n2;
	CLB_3_2_IN_pin_4_driver_mux_fanins <= track_3_2_chanX_n11 & track_3_2_chanX_n10 & track_3_2_chanX_n3 & track_3_2_chanX_n2;
	CLB_3_2_IN_pin_5_driver_mux_fanins <= track_3_2_chanY_n13 & track_3_2_chanY_n12 & track_3_2_chanY_n5 & track_3_2_chanY_n4;
	CLB_3_2_IN_pin_6_driver_mux_fanins <= track_3_1_chanX_n13 & track_3_1_chanX_n12 & track_3_1_chanX_n5 & track_3_1_chanX_n4;
	CLB_3_2_IN_pin_7_driver_mux_fanins <= track_2_2_chanY_n13 & track_2_2_chanY_n12 & track_2_2_chanY_n5 & track_2_2_chanY_n4;
	CLB_3_2_IN_pin_8_driver_mux_fanins <= track_3_2_chanX_n15 & track_3_2_chanX_n14 & track_3_2_chanX_n7 & track_3_2_chanX_n6;
	CLB_3_2_IN_pin_9_driver_mux_fanins <= track_3_2_chanY_n15 & track_3_2_chanY_n14 & track_3_2_chanY_n7 & track_3_2_chanY_n6;
	CLB_3_3_IN_pin_0_driver_mux_fanins <= track_3_3_chanX_n9 & track_3_3_chanX_n8 & track_3_3_chanX_n1 & track_3_3_chanX_n0;
	CLB_3_3_IN_pin_1_driver_mux_fanins <= track_3_3_chanY_n9 & track_3_3_chanY_n8 & track_3_3_chanY_n1 & track_3_3_chanY_n0;
	CLB_3_3_IN_pin_2_driver_mux_fanins <= track_3_2_chanX_n9 & track_3_2_chanX_n8 & track_3_2_chanX_n1 & track_3_2_chanX_n0;
	CLB_3_3_IN_pin_3_driver_mux_fanins <= track_2_3_chanY_n11 & track_2_3_chanY_n10 & track_2_3_chanY_n3 & track_2_3_chanY_n2;
	CLB_3_3_IN_pin_4_driver_mux_fanins <= track_3_3_chanX_n11 & track_3_3_chanX_n10 & track_3_3_chanX_n3 & track_3_3_chanX_n2;
	CLB_3_3_IN_pin_5_driver_mux_fanins <= track_3_3_chanY_n13 & track_3_3_chanY_n12 & track_3_3_chanY_n5 & track_3_3_chanY_n4;
	CLB_3_3_IN_pin_6_driver_mux_fanins <= track_3_2_chanX_n13 & track_3_2_chanX_n12 & track_3_2_chanX_n5 & track_3_2_chanX_n4;
	CLB_3_3_IN_pin_7_driver_mux_fanins <= track_2_3_chanY_n13 & track_2_3_chanY_n12 & track_2_3_chanY_n5 & track_2_3_chanY_n4;
	CLB_3_3_IN_pin_8_driver_mux_fanins <= track_3_3_chanX_n15 & track_3_3_chanX_n14 & track_3_3_chanX_n7 & track_3_3_chanX_n6;
	CLB_3_3_IN_pin_9_driver_mux_fanins <= track_3_3_chanY_n15 & track_3_3_chanY_n14 & track_3_3_chanY_n7 & track_3_3_chanY_n6;
	CLB_3_4_IN_pin_0_driver_mux_fanins <= track_3_4_chanX_n9 & track_3_4_chanX_n8 & track_3_4_chanX_n1 & track_3_4_chanX_n0;
	CLB_3_4_IN_pin_1_driver_mux_fanins <= track_3_4_chanY_n9 & track_3_4_chanY_n8 & track_3_4_chanY_n1 & track_3_4_chanY_n0;
	CLB_3_4_IN_pin_2_driver_mux_fanins <= track_3_3_chanX_n9 & track_3_3_chanX_n8 & track_3_3_chanX_n1 & track_3_3_chanX_n0;
	CLB_3_4_IN_pin_3_driver_mux_fanins <= track_2_4_chanY_n11 & track_2_4_chanY_n10 & track_2_4_chanY_n3 & track_2_4_chanY_n2;
	CLB_3_4_IN_pin_4_driver_mux_fanins <= track_3_4_chanX_n11 & track_3_4_chanX_n10 & track_3_4_chanX_n3 & track_3_4_chanX_n2;
	CLB_3_4_IN_pin_5_driver_mux_fanins <= track_3_4_chanY_n13 & track_3_4_chanY_n12 & track_3_4_chanY_n5 & track_3_4_chanY_n4;
	CLB_3_4_IN_pin_6_driver_mux_fanins <= track_3_3_chanX_n13 & track_3_3_chanX_n12 & track_3_3_chanX_n5 & track_3_3_chanX_n4;
	CLB_3_4_IN_pin_7_driver_mux_fanins <= track_2_4_chanY_n13 & track_2_4_chanY_n12 & track_2_4_chanY_n5 & track_2_4_chanY_n4;
	CLB_3_4_IN_pin_8_driver_mux_fanins <= track_3_4_chanX_n15 & track_3_4_chanX_n14 & track_3_4_chanX_n7 & track_3_4_chanX_n6;
	CLB_3_4_IN_pin_9_driver_mux_fanins <= track_3_4_chanY_n15 & track_3_4_chanY_n14 & track_3_4_chanY_n7 & track_3_4_chanY_n6;
	CLB_3_5_IN_pin_0_driver_mux_fanins <= track_3_5_chanX_n9 & track_3_5_chanX_n8 & track_3_5_chanX_n1 & track_3_5_chanX_n0;
	CLB_3_5_IN_pin_1_driver_mux_fanins <= track_3_5_chanY_n9 & track_3_5_chanY_n8 & track_3_5_chanY_n1 & track_3_5_chanY_n0;
	CLB_3_5_IN_pin_2_driver_mux_fanins <= track_3_4_chanX_n9 & track_3_4_chanX_n8 & track_3_4_chanX_n1 & track_3_4_chanX_n0;
	CLB_3_5_IN_pin_3_driver_mux_fanins <= track_2_5_chanY_n11 & track_2_5_chanY_n10 & track_2_5_chanY_n3 & track_2_5_chanY_n2;
	CLB_3_5_IN_pin_4_driver_mux_fanins <= track_3_5_chanX_n11 & track_3_5_chanX_n10 & track_3_5_chanX_n3 & track_3_5_chanX_n2;
	CLB_3_5_IN_pin_5_driver_mux_fanins <= track_3_5_chanY_n13 & track_3_5_chanY_n12 & track_3_5_chanY_n5 & track_3_5_chanY_n4;
	CLB_3_5_IN_pin_6_driver_mux_fanins <= track_3_4_chanX_n13 & track_3_4_chanX_n12 & track_3_4_chanX_n5 & track_3_4_chanX_n4;
	CLB_3_5_IN_pin_7_driver_mux_fanins <= track_2_5_chanY_n13 & track_2_5_chanY_n12 & track_2_5_chanY_n5 & track_2_5_chanY_n4;
	CLB_3_5_IN_pin_8_driver_mux_fanins <= track_3_5_chanX_n15 & track_3_5_chanX_n14 & track_3_5_chanX_n7 & track_3_5_chanX_n6;
	CLB_3_5_IN_pin_9_driver_mux_fanins <= track_3_5_chanY_n15 & track_3_5_chanY_n14 & track_3_5_chanY_n7 & track_3_5_chanY_n6;
	CLB_3_6_IN_pin_0_driver_mux_fanins <= track_3_6_chanX_n9 & track_3_6_chanX_n8 & track_3_6_chanX_n1 & track_3_6_chanX_n0;
	CLB_3_6_IN_pin_1_driver_mux_fanins <= track_3_6_chanY_n9 & track_3_6_chanY_n8 & track_3_6_chanY_n1 & track_3_6_chanY_n0;
	CLB_3_6_IN_pin_2_driver_mux_fanins <= track_3_5_chanX_n9 & track_3_5_chanX_n8 & track_3_5_chanX_n1 & track_3_5_chanX_n0;
	CLB_3_6_IN_pin_3_driver_mux_fanins <= track_2_6_chanY_n11 & track_2_6_chanY_n10 & track_2_6_chanY_n3 & track_2_6_chanY_n2;
	CLB_3_6_IN_pin_4_driver_mux_fanins <= track_3_6_chanX_n11 & track_3_6_chanX_n10 & track_3_6_chanX_n3 & track_3_6_chanX_n2;
	CLB_3_6_IN_pin_5_driver_mux_fanins <= track_3_6_chanY_n13 & track_3_6_chanY_n12 & track_3_6_chanY_n5 & track_3_6_chanY_n4;
	CLB_3_6_IN_pin_6_driver_mux_fanins <= track_3_5_chanX_n13 & track_3_5_chanX_n12 & track_3_5_chanX_n5 & track_3_5_chanX_n4;
	CLB_3_6_IN_pin_7_driver_mux_fanins <= track_2_6_chanY_n13 & track_2_6_chanY_n12 & track_2_6_chanY_n5 & track_2_6_chanY_n4;
	CLB_3_6_IN_pin_8_driver_mux_fanins <= track_3_6_chanX_n15 & track_3_6_chanX_n14 & track_3_6_chanX_n7 & track_3_6_chanX_n6;
	CLB_3_6_IN_pin_9_driver_mux_fanins <= track_3_6_chanY_n15 & track_3_6_chanY_n14 & track_3_6_chanY_n7 & track_3_6_chanY_n6;
	CLB_4_1_IN_pin_0_driver_mux_fanins <= track_4_1_chanX_n9 & track_4_1_chanX_n8 & track_4_1_chanX_n1 & track_4_1_chanX_n0;
	CLB_4_1_IN_pin_1_driver_mux_fanins <= track_4_1_chanY_n9 & track_4_1_chanY_n8 & track_4_1_chanY_n1 & track_4_1_chanY_n0;
	CLB_4_1_IN_pin_2_driver_mux_fanins <= track_4_0_chanX_n9 & track_4_0_chanX_n8 & track_4_0_chanX_n1 & track_4_0_chanX_n0;
	CLB_4_1_IN_pin_3_driver_mux_fanins <= track_3_1_chanY_n11 & track_3_1_chanY_n10 & track_3_1_chanY_n3 & track_3_1_chanY_n2;
	CLB_4_1_IN_pin_4_driver_mux_fanins <= track_4_1_chanX_n11 & track_4_1_chanX_n10 & track_4_1_chanX_n3 & track_4_1_chanX_n2;
	CLB_4_1_IN_pin_5_driver_mux_fanins <= track_4_1_chanY_n13 & track_4_1_chanY_n12 & track_4_1_chanY_n5 & track_4_1_chanY_n4;
	CLB_4_1_IN_pin_6_driver_mux_fanins <= track_4_0_chanX_n13 & track_4_0_chanX_n12 & track_4_0_chanX_n5 & track_4_0_chanX_n4;
	CLB_4_1_IN_pin_7_driver_mux_fanins <= track_3_1_chanY_n13 & track_3_1_chanY_n12 & track_3_1_chanY_n5 & track_3_1_chanY_n4;
	CLB_4_1_IN_pin_8_driver_mux_fanins <= track_4_1_chanX_n15 & track_4_1_chanX_n14 & track_4_1_chanX_n7 & track_4_1_chanX_n6;
	CLB_4_1_IN_pin_9_driver_mux_fanins <= track_4_1_chanY_n15 & track_4_1_chanY_n14 & track_4_1_chanY_n7 & track_4_1_chanY_n6;
	CLB_4_2_IN_pin_0_driver_mux_fanins <= track_4_2_chanX_n9 & track_4_2_chanX_n8 & track_4_2_chanX_n1 & track_4_2_chanX_n0;
	CLB_4_2_IN_pin_1_driver_mux_fanins <= track_4_2_chanY_n9 & track_4_2_chanY_n8 & track_4_2_chanY_n1 & track_4_2_chanY_n0;
	CLB_4_2_IN_pin_2_driver_mux_fanins <= track_4_1_chanX_n9 & track_4_1_chanX_n8 & track_4_1_chanX_n1 & track_4_1_chanX_n0;
	CLB_4_2_IN_pin_3_driver_mux_fanins <= track_3_2_chanY_n11 & track_3_2_chanY_n10 & track_3_2_chanY_n3 & track_3_2_chanY_n2;
	CLB_4_2_IN_pin_4_driver_mux_fanins <= track_4_2_chanX_n11 & track_4_2_chanX_n10 & track_4_2_chanX_n3 & track_4_2_chanX_n2;
	CLB_4_2_IN_pin_5_driver_mux_fanins <= track_4_2_chanY_n13 & track_4_2_chanY_n12 & track_4_2_chanY_n5 & track_4_2_chanY_n4;
	CLB_4_2_IN_pin_6_driver_mux_fanins <= track_4_1_chanX_n13 & track_4_1_chanX_n12 & track_4_1_chanX_n5 & track_4_1_chanX_n4;
	CLB_4_2_IN_pin_7_driver_mux_fanins <= track_3_2_chanY_n13 & track_3_2_chanY_n12 & track_3_2_chanY_n5 & track_3_2_chanY_n4;
	CLB_4_2_IN_pin_8_driver_mux_fanins <= track_4_2_chanX_n15 & track_4_2_chanX_n14 & track_4_2_chanX_n7 & track_4_2_chanX_n6;
	CLB_4_2_IN_pin_9_driver_mux_fanins <= track_4_2_chanY_n15 & track_4_2_chanY_n14 & track_4_2_chanY_n7 & track_4_2_chanY_n6;
	CLB_4_3_IN_pin_0_driver_mux_fanins <= track_4_3_chanX_n9 & track_4_3_chanX_n8 & track_4_3_chanX_n1 & track_4_3_chanX_n0;
	CLB_4_3_IN_pin_1_driver_mux_fanins <= track_4_3_chanY_n9 & track_4_3_chanY_n8 & track_4_3_chanY_n1 & track_4_3_chanY_n0;
	CLB_4_3_IN_pin_2_driver_mux_fanins <= track_4_2_chanX_n9 & track_4_2_chanX_n8 & track_4_2_chanX_n1 & track_4_2_chanX_n0;
	CLB_4_3_IN_pin_3_driver_mux_fanins <= track_3_3_chanY_n11 & track_3_3_chanY_n10 & track_3_3_chanY_n3 & track_3_3_chanY_n2;
	CLB_4_3_IN_pin_4_driver_mux_fanins <= track_4_3_chanX_n11 & track_4_3_chanX_n10 & track_4_3_chanX_n3 & track_4_3_chanX_n2;
	CLB_4_3_IN_pin_5_driver_mux_fanins <= track_4_3_chanY_n13 & track_4_3_chanY_n12 & track_4_3_chanY_n5 & track_4_3_chanY_n4;
	CLB_4_3_IN_pin_6_driver_mux_fanins <= track_4_2_chanX_n13 & track_4_2_chanX_n12 & track_4_2_chanX_n5 & track_4_2_chanX_n4;
	CLB_4_3_IN_pin_7_driver_mux_fanins <= track_3_3_chanY_n13 & track_3_3_chanY_n12 & track_3_3_chanY_n5 & track_3_3_chanY_n4;
	CLB_4_3_IN_pin_8_driver_mux_fanins <= track_4_3_chanX_n15 & track_4_3_chanX_n14 & track_4_3_chanX_n7 & track_4_3_chanX_n6;
	CLB_4_3_IN_pin_9_driver_mux_fanins <= track_4_3_chanY_n15 & track_4_3_chanY_n14 & track_4_3_chanY_n7 & track_4_3_chanY_n6;
	CLB_4_4_IN_pin_0_driver_mux_fanins <= track_4_4_chanX_n9 & track_4_4_chanX_n8 & track_4_4_chanX_n1 & track_4_4_chanX_n0;
	CLB_4_4_IN_pin_1_driver_mux_fanins <= track_4_4_chanY_n9 & track_4_4_chanY_n8 & track_4_4_chanY_n1 & track_4_4_chanY_n0;
	CLB_4_4_IN_pin_2_driver_mux_fanins <= track_4_3_chanX_n9 & track_4_3_chanX_n8 & track_4_3_chanX_n1 & track_4_3_chanX_n0;
	CLB_4_4_IN_pin_3_driver_mux_fanins <= track_3_4_chanY_n11 & track_3_4_chanY_n10 & track_3_4_chanY_n3 & track_3_4_chanY_n2;
	CLB_4_4_IN_pin_4_driver_mux_fanins <= track_4_4_chanX_n11 & track_4_4_chanX_n10 & track_4_4_chanX_n3 & track_4_4_chanX_n2;
	CLB_4_4_IN_pin_5_driver_mux_fanins <= track_4_4_chanY_n13 & track_4_4_chanY_n12 & track_4_4_chanY_n5 & track_4_4_chanY_n4;
	CLB_4_4_IN_pin_6_driver_mux_fanins <= track_4_3_chanX_n13 & track_4_3_chanX_n12 & track_4_3_chanX_n5 & track_4_3_chanX_n4;
	CLB_4_4_IN_pin_7_driver_mux_fanins <= track_3_4_chanY_n13 & track_3_4_chanY_n12 & track_3_4_chanY_n5 & track_3_4_chanY_n4;
	CLB_4_4_IN_pin_8_driver_mux_fanins <= track_4_4_chanX_n15 & track_4_4_chanX_n14 & track_4_4_chanX_n7 & track_4_4_chanX_n6;
	CLB_4_4_IN_pin_9_driver_mux_fanins <= track_4_4_chanY_n15 & track_4_4_chanY_n14 & track_4_4_chanY_n7 & track_4_4_chanY_n6;
	CLB_4_5_IN_pin_0_driver_mux_fanins <= track_4_5_chanX_n9 & track_4_5_chanX_n8 & track_4_5_chanX_n1 & track_4_5_chanX_n0;
	CLB_4_5_IN_pin_1_driver_mux_fanins <= track_4_5_chanY_n9 & track_4_5_chanY_n8 & track_4_5_chanY_n1 & track_4_5_chanY_n0;
	CLB_4_5_IN_pin_2_driver_mux_fanins <= track_4_4_chanX_n9 & track_4_4_chanX_n8 & track_4_4_chanX_n1 & track_4_4_chanX_n0;
	CLB_4_5_IN_pin_3_driver_mux_fanins <= track_3_5_chanY_n11 & track_3_5_chanY_n10 & track_3_5_chanY_n3 & track_3_5_chanY_n2;
	CLB_4_5_IN_pin_4_driver_mux_fanins <= track_4_5_chanX_n11 & track_4_5_chanX_n10 & track_4_5_chanX_n3 & track_4_5_chanX_n2;
	CLB_4_5_IN_pin_5_driver_mux_fanins <= track_4_5_chanY_n13 & track_4_5_chanY_n12 & track_4_5_chanY_n5 & track_4_5_chanY_n4;
	CLB_4_5_IN_pin_6_driver_mux_fanins <= track_4_4_chanX_n13 & track_4_4_chanX_n12 & track_4_4_chanX_n5 & track_4_4_chanX_n4;
	CLB_4_5_IN_pin_7_driver_mux_fanins <= track_3_5_chanY_n13 & track_3_5_chanY_n12 & track_3_5_chanY_n5 & track_3_5_chanY_n4;
	CLB_4_5_IN_pin_8_driver_mux_fanins <= track_4_5_chanX_n15 & track_4_5_chanX_n14 & track_4_5_chanX_n7 & track_4_5_chanX_n6;
	CLB_4_5_IN_pin_9_driver_mux_fanins <= track_4_5_chanY_n15 & track_4_5_chanY_n14 & track_4_5_chanY_n7 & track_4_5_chanY_n6;
	CLB_4_6_IN_pin_0_driver_mux_fanins <= track_4_6_chanX_n9 & track_4_6_chanX_n8 & track_4_6_chanX_n1 & track_4_6_chanX_n0;
	CLB_4_6_IN_pin_1_driver_mux_fanins <= track_4_6_chanY_n9 & track_4_6_chanY_n8 & track_4_6_chanY_n1 & track_4_6_chanY_n0;
	CLB_4_6_IN_pin_2_driver_mux_fanins <= track_4_5_chanX_n9 & track_4_5_chanX_n8 & track_4_5_chanX_n1 & track_4_5_chanX_n0;
	CLB_4_6_IN_pin_3_driver_mux_fanins <= track_3_6_chanY_n11 & track_3_6_chanY_n10 & track_3_6_chanY_n3 & track_3_6_chanY_n2;
	CLB_4_6_IN_pin_4_driver_mux_fanins <= track_4_6_chanX_n11 & track_4_6_chanX_n10 & track_4_6_chanX_n3 & track_4_6_chanX_n2;
	CLB_4_6_IN_pin_5_driver_mux_fanins <= track_4_6_chanY_n13 & track_4_6_chanY_n12 & track_4_6_chanY_n5 & track_4_6_chanY_n4;
	CLB_4_6_IN_pin_6_driver_mux_fanins <= track_4_5_chanX_n13 & track_4_5_chanX_n12 & track_4_5_chanX_n5 & track_4_5_chanX_n4;
	CLB_4_6_IN_pin_7_driver_mux_fanins <= track_3_6_chanY_n13 & track_3_6_chanY_n12 & track_3_6_chanY_n5 & track_3_6_chanY_n4;
	CLB_4_6_IN_pin_8_driver_mux_fanins <= track_4_6_chanX_n15 & track_4_6_chanX_n14 & track_4_6_chanX_n7 & track_4_6_chanX_n6;
	CLB_4_6_IN_pin_9_driver_mux_fanins <= track_4_6_chanY_n15 & track_4_6_chanY_n14 & track_4_6_chanY_n7 & track_4_6_chanY_n6;
	CLB_5_1_IN_pin_0_driver_mux_fanins <= track_5_1_chanX_n9 & track_5_1_chanX_n8 & track_5_1_chanX_n1 & track_5_1_chanX_n0;
	CLB_5_1_IN_pin_1_driver_mux_fanins <= track_5_1_chanY_n9 & track_5_1_chanY_n8 & track_5_1_chanY_n1 & track_5_1_chanY_n0;
	CLB_5_1_IN_pin_2_driver_mux_fanins <= track_5_0_chanX_n9 & track_5_0_chanX_n8 & track_5_0_chanX_n1 & track_5_0_chanX_n0;
	CLB_5_1_IN_pin_3_driver_mux_fanins <= track_4_1_chanY_n11 & track_4_1_chanY_n10 & track_4_1_chanY_n3 & track_4_1_chanY_n2;
	CLB_5_1_IN_pin_4_driver_mux_fanins <= track_5_1_chanX_n11 & track_5_1_chanX_n10 & track_5_1_chanX_n3 & track_5_1_chanX_n2;
	CLB_5_1_IN_pin_5_driver_mux_fanins <= track_5_1_chanY_n13 & track_5_1_chanY_n12 & track_5_1_chanY_n5 & track_5_1_chanY_n4;
	CLB_5_1_IN_pin_6_driver_mux_fanins <= track_5_0_chanX_n13 & track_5_0_chanX_n12 & track_5_0_chanX_n5 & track_5_0_chanX_n4;
	CLB_5_1_IN_pin_7_driver_mux_fanins <= track_4_1_chanY_n13 & track_4_1_chanY_n12 & track_4_1_chanY_n5 & track_4_1_chanY_n4;
	CLB_5_1_IN_pin_8_driver_mux_fanins <= track_5_1_chanX_n15 & track_5_1_chanX_n14 & track_5_1_chanX_n7 & track_5_1_chanX_n6;
	CLB_5_1_IN_pin_9_driver_mux_fanins <= track_5_1_chanY_n15 & track_5_1_chanY_n14 & track_5_1_chanY_n7 & track_5_1_chanY_n6;
	CLB_5_2_IN_pin_0_driver_mux_fanins <= track_5_2_chanX_n9 & track_5_2_chanX_n8 & track_5_2_chanX_n1 & track_5_2_chanX_n0;
	CLB_5_2_IN_pin_1_driver_mux_fanins <= track_5_2_chanY_n9 & track_5_2_chanY_n8 & track_5_2_chanY_n1 & track_5_2_chanY_n0;
	CLB_5_2_IN_pin_2_driver_mux_fanins <= track_5_1_chanX_n9 & track_5_1_chanX_n8 & track_5_1_chanX_n1 & track_5_1_chanX_n0;
	CLB_5_2_IN_pin_3_driver_mux_fanins <= track_4_2_chanY_n11 & track_4_2_chanY_n10 & track_4_2_chanY_n3 & track_4_2_chanY_n2;
	CLB_5_2_IN_pin_4_driver_mux_fanins <= track_5_2_chanX_n11 & track_5_2_chanX_n10 & track_5_2_chanX_n3 & track_5_2_chanX_n2;
	CLB_5_2_IN_pin_5_driver_mux_fanins <= track_5_2_chanY_n13 & track_5_2_chanY_n12 & track_5_2_chanY_n5 & track_5_2_chanY_n4;
	CLB_5_2_IN_pin_6_driver_mux_fanins <= track_5_1_chanX_n13 & track_5_1_chanX_n12 & track_5_1_chanX_n5 & track_5_1_chanX_n4;
	CLB_5_2_IN_pin_7_driver_mux_fanins <= track_4_2_chanY_n13 & track_4_2_chanY_n12 & track_4_2_chanY_n5 & track_4_2_chanY_n4;
	CLB_5_2_IN_pin_8_driver_mux_fanins <= track_5_2_chanX_n15 & track_5_2_chanX_n14 & track_5_2_chanX_n7 & track_5_2_chanX_n6;
	CLB_5_2_IN_pin_9_driver_mux_fanins <= track_5_2_chanY_n15 & track_5_2_chanY_n14 & track_5_2_chanY_n7 & track_5_2_chanY_n6;
	CLB_5_3_IN_pin_0_driver_mux_fanins <= track_5_3_chanX_n9 & track_5_3_chanX_n8 & track_5_3_chanX_n1 & track_5_3_chanX_n0;
	CLB_5_3_IN_pin_1_driver_mux_fanins <= track_5_3_chanY_n9 & track_5_3_chanY_n8 & track_5_3_chanY_n1 & track_5_3_chanY_n0;
	CLB_5_3_IN_pin_2_driver_mux_fanins <= track_5_2_chanX_n9 & track_5_2_chanX_n8 & track_5_2_chanX_n1 & track_5_2_chanX_n0;
	CLB_5_3_IN_pin_3_driver_mux_fanins <= track_4_3_chanY_n11 & track_4_3_chanY_n10 & track_4_3_chanY_n3 & track_4_3_chanY_n2;
	CLB_5_3_IN_pin_4_driver_mux_fanins <= track_5_3_chanX_n11 & track_5_3_chanX_n10 & track_5_3_chanX_n3 & track_5_3_chanX_n2;
	CLB_5_3_IN_pin_5_driver_mux_fanins <= track_5_3_chanY_n13 & track_5_3_chanY_n12 & track_5_3_chanY_n5 & track_5_3_chanY_n4;
	CLB_5_3_IN_pin_6_driver_mux_fanins <= track_5_2_chanX_n13 & track_5_2_chanX_n12 & track_5_2_chanX_n5 & track_5_2_chanX_n4;
	CLB_5_3_IN_pin_7_driver_mux_fanins <= track_4_3_chanY_n13 & track_4_3_chanY_n12 & track_4_3_chanY_n5 & track_4_3_chanY_n4;
	CLB_5_3_IN_pin_8_driver_mux_fanins <= track_5_3_chanX_n15 & track_5_3_chanX_n14 & track_5_3_chanX_n7 & track_5_3_chanX_n6;
	CLB_5_3_IN_pin_9_driver_mux_fanins <= track_5_3_chanY_n15 & track_5_3_chanY_n14 & track_5_3_chanY_n7 & track_5_3_chanY_n6;
	CLB_5_4_IN_pin_0_driver_mux_fanins <= track_5_4_chanX_n9 & track_5_4_chanX_n8 & track_5_4_chanX_n1 & track_5_4_chanX_n0;
	CLB_5_4_IN_pin_1_driver_mux_fanins <= track_5_4_chanY_n9 & track_5_4_chanY_n8 & track_5_4_chanY_n1 & track_5_4_chanY_n0;
	CLB_5_4_IN_pin_2_driver_mux_fanins <= track_5_3_chanX_n9 & track_5_3_chanX_n8 & track_5_3_chanX_n1 & track_5_3_chanX_n0;
	CLB_5_4_IN_pin_3_driver_mux_fanins <= track_4_4_chanY_n11 & track_4_4_chanY_n10 & track_4_4_chanY_n3 & track_4_4_chanY_n2;
	CLB_5_4_IN_pin_4_driver_mux_fanins <= track_5_4_chanX_n11 & track_5_4_chanX_n10 & track_5_4_chanX_n3 & track_5_4_chanX_n2;
	CLB_5_4_IN_pin_5_driver_mux_fanins <= track_5_4_chanY_n13 & track_5_4_chanY_n12 & track_5_4_chanY_n5 & track_5_4_chanY_n4;
	CLB_5_4_IN_pin_6_driver_mux_fanins <= track_5_3_chanX_n13 & track_5_3_chanX_n12 & track_5_3_chanX_n5 & track_5_3_chanX_n4;
	CLB_5_4_IN_pin_7_driver_mux_fanins <= track_4_4_chanY_n13 & track_4_4_chanY_n12 & track_4_4_chanY_n5 & track_4_4_chanY_n4;
	CLB_5_4_IN_pin_8_driver_mux_fanins <= track_5_4_chanX_n15 & track_5_4_chanX_n14 & track_5_4_chanX_n7 & track_5_4_chanX_n6;
	CLB_5_4_IN_pin_9_driver_mux_fanins <= track_5_4_chanY_n15 & track_5_4_chanY_n14 & track_5_4_chanY_n7 & track_5_4_chanY_n6;
	CLB_5_5_IN_pin_0_driver_mux_fanins <= track_5_5_chanX_n9 & track_5_5_chanX_n8 & track_5_5_chanX_n1 & track_5_5_chanX_n0;
	CLB_5_5_IN_pin_1_driver_mux_fanins <= track_5_5_chanY_n9 & track_5_5_chanY_n8 & track_5_5_chanY_n1 & track_5_5_chanY_n0;
	CLB_5_5_IN_pin_2_driver_mux_fanins <= track_5_4_chanX_n9 & track_5_4_chanX_n8 & track_5_4_chanX_n1 & track_5_4_chanX_n0;
	CLB_5_5_IN_pin_3_driver_mux_fanins <= track_4_5_chanY_n11 & track_4_5_chanY_n10 & track_4_5_chanY_n3 & track_4_5_chanY_n2;
	CLB_5_5_IN_pin_4_driver_mux_fanins <= track_5_5_chanX_n11 & track_5_5_chanX_n10 & track_5_5_chanX_n3 & track_5_5_chanX_n2;
	CLB_5_5_IN_pin_5_driver_mux_fanins <= track_5_5_chanY_n13 & track_5_5_chanY_n12 & track_5_5_chanY_n5 & track_5_5_chanY_n4;
	CLB_5_5_IN_pin_6_driver_mux_fanins <= track_5_4_chanX_n13 & track_5_4_chanX_n12 & track_5_4_chanX_n5 & track_5_4_chanX_n4;
	CLB_5_5_IN_pin_7_driver_mux_fanins <= track_4_5_chanY_n13 & track_4_5_chanY_n12 & track_4_5_chanY_n5 & track_4_5_chanY_n4;
	CLB_5_5_IN_pin_8_driver_mux_fanins <= track_5_5_chanX_n15 & track_5_5_chanX_n14 & track_5_5_chanX_n7 & track_5_5_chanX_n6;
	CLB_5_5_IN_pin_9_driver_mux_fanins <= track_5_5_chanY_n15 & track_5_5_chanY_n14 & track_5_5_chanY_n7 & track_5_5_chanY_n6;
	CLB_5_6_IN_pin_0_driver_mux_fanins <= track_5_6_chanX_n9 & track_5_6_chanX_n8 & track_5_6_chanX_n1 & track_5_6_chanX_n0;
	CLB_5_6_IN_pin_1_driver_mux_fanins <= track_5_6_chanY_n9 & track_5_6_chanY_n8 & track_5_6_chanY_n1 & track_5_6_chanY_n0;
	CLB_5_6_IN_pin_2_driver_mux_fanins <= track_5_5_chanX_n9 & track_5_5_chanX_n8 & track_5_5_chanX_n1 & track_5_5_chanX_n0;
	CLB_5_6_IN_pin_3_driver_mux_fanins <= track_4_6_chanY_n11 & track_4_6_chanY_n10 & track_4_6_chanY_n3 & track_4_6_chanY_n2;
	CLB_5_6_IN_pin_4_driver_mux_fanins <= track_5_6_chanX_n11 & track_5_6_chanX_n10 & track_5_6_chanX_n3 & track_5_6_chanX_n2;
	CLB_5_6_IN_pin_5_driver_mux_fanins <= track_5_6_chanY_n13 & track_5_6_chanY_n12 & track_5_6_chanY_n5 & track_5_6_chanY_n4;
	CLB_5_6_IN_pin_6_driver_mux_fanins <= track_5_5_chanX_n13 & track_5_5_chanX_n12 & track_5_5_chanX_n5 & track_5_5_chanX_n4;
	CLB_5_6_IN_pin_7_driver_mux_fanins <= track_4_6_chanY_n13 & track_4_6_chanY_n12 & track_4_6_chanY_n5 & track_4_6_chanY_n4;
	CLB_5_6_IN_pin_8_driver_mux_fanins <= track_5_6_chanX_n15 & track_5_6_chanX_n14 & track_5_6_chanX_n7 & track_5_6_chanX_n6;
	CLB_5_6_IN_pin_9_driver_mux_fanins <= track_5_6_chanY_n15 & track_5_6_chanY_n14 & track_5_6_chanY_n7 & track_5_6_chanY_n6;
	CLB_6_1_IN_pin_0_driver_mux_fanins <= track_6_1_chanX_n9 & track_6_1_chanX_n8 & track_6_1_chanX_n1 & track_6_1_chanX_n0;
	CLB_6_1_IN_pin_1_driver_mux_fanins <= track_6_1_chanY_n9 & track_6_1_chanY_n8 & track_6_1_chanY_n1 & track_6_1_chanY_n0;
	CLB_6_1_IN_pin_2_driver_mux_fanins <= track_6_0_chanX_n9 & track_6_0_chanX_n8 & track_6_0_chanX_n1 & track_6_0_chanX_n0;
	CLB_6_1_IN_pin_3_driver_mux_fanins <= track_5_1_chanY_n11 & track_5_1_chanY_n10 & track_5_1_chanY_n3 & track_5_1_chanY_n2;
	CLB_6_1_IN_pin_4_driver_mux_fanins <= track_6_1_chanX_n11 & track_6_1_chanX_n10 & track_6_1_chanX_n3 & track_6_1_chanX_n2;
	CLB_6_1_IN_pin_5_driver_mux_fanins <= track_6_1_chanY_n13 & track_6_1_chanY_n12 & track_6_1_chanY_n5 & track_6_1_chanY_n4;
	CLB_6_1_IN_pin_6_driver_mux_fanins <= track_6_0_chanX_n13 & track_6_0_chanX_n12 & track_6_0_chanX_n5 & track_6_0_chanX_n4;
	CLB_6_1_IN_pin_7_driver_mux_fanins <= track_5_1_chanY_n13 & track_5_1_chanY_n12 & track_5_1_chanY_n5 & track_5_1_chanY_n4;
	CLB_6_1_IN_pin_8_driver_mux_fanins <= track_6_1_chanX_n15 & track_6_1_chanX_n14 & track_6_1_chanX_n7 & track_6_1_chanX_n6;
	CLB_6_1_IN_pin_9_driver_mux_fanins <= track_6_1_chanY_n15 & track_6_1_chanY_n14 & track_6_1_chanY_n7 & track_6_1_chanY_n6;
	CLB_6_2_IN_pin_0_driver_mux_fanins <= track_6_2_chanX_n9 & track_6_2_chanX_n8 & track_6_2_chanX_n1 & track_6_2_chanX_n0;
	CLB_6_2_IN_pin_1_driver_mux_fanins <= track_6_2_chanY_n9 & track_6_2_chanY_n8 & track_6_2_chanY_n1 & track_6_2_chanY_n0;
	CLB_6_2_IN_pin_2_driver_mux_fanins <= track_6_1_chanX_n9 & track_6_1_chanX_n8 & track_6_1_chanX_n1 & track_6_1_chanX_n0;
	CLB_6_2_IN_pin_3_driver_mux_fanins <= track_5_2_chanY_n11 & track_5_2_chanY_n10 & track_5_2_chanY_n3 & track_5_2_chanY_n2;
	CLB_6_2_IN_pin_4_driver_mux_fanins <= track_6_2_chanX_n11 & track_6_2_chanX_n10 & track_6_2_chanX_n3 & track_6_2_chanX_n2;
	CLB_6_2_IN_pin_5_driver_mux_fanins <= track_6_2_chanY_n13 & track_6_2_chanY_n12 & track_6_2_chanY_n5 & track_6_2_chanY_n4;
	CLB_6_2_IN_pin_6_driver_mux_fanins <= track_6_1_chanX_n13 & track_6_1_chanX_n12 & track_6_1_chanX_n5 & track_6_1_chanX_n4;
	CLB_6_2_IN_pin_7_driver_mux_fanins <= track_5_2_chanY_n13 & track_5_2_chanY_n12 & track_5_2_chanY_n5 & track_5_2_chanY_n4;
	CLB_6_2_IN_pin_8_driver_mux_fanins <= track_6_2_chanX_n15 & track_6_2_chanX_n14 & track_6_2_chanX_n7 & track_6_2_chanX_n6;
	CLB_6_2_IN_pin_9_driver_mux_fanins <= track_6_2_chanY_n15 & track_6_2_chanY_n14 & track_6_2_chanY_n7 & track_6_2_chanY_n6;
	CLB_6_3_IN_pin_0_driver_mux_fanins <= track_6_3_chanX_n9 & track_6_3_chanX_n8 & track_6_3_chanX_n1 & track_6_3_chanX_n0;
	CLB_6_3_IN_pin_1_driver_mux_fanins <= track_6_3_chanY_n9 & track_6_3_chanY_n8 & track_6_3_chanY_n1 & track_6_3_chanY_n0;
	CLB_6_3_IN_pin_2_driver_mux_fanins <= track_6_2_chanX_n9 & track_6_2_chanX_n8 & track_6_2_chanX_n1 & track_6_2_chanX_n0;
	CLB_6_3_IN_pin_3_driver_mux_fanins <= track_5_3_chanY_n11 & track_5_3_chanY_n10 & track_5_3_chanY_n3 & track_5_3_chanY_n2;
	CLB_6_3_IN_pin_4_driver_mux_fanins <= track_6_3_chanX_n11 & track_6_3_chanX_n10 & track_6_3_chanX_n3 & track_6_3_chanX_n2;
	CLB_6_3_IN_pin_5_driver_mux_fanins <= track_6_3_chanY_n13 & track_6_3_chanY_n12 & track_6_3_chanY_n5 & track_6_3_chanY_n4;
	CLB_6_3_IN_pin_6_driver_mux_fanins <= track_6_2_chanX_n13 & track_6_2_chanX_n12 & track_6_2_chanX_n5 & track_6_2_chanX_n4;
	CLB_6_3_IN_pin_7_driver_mux_fanins <= track_5_3_chanY_n13 & track_5_3_chanY_n12 & track_5_3_chanY_n5 & track_5_3_chanY_n4;
	CLB_6_3_IN_pin_8_driver_mux_fanins <= track_6_3_chanX_n15 & track_6_3_chanX_n14 & track_6_3_chanX_n7 & track_6_3_chanX_n6;
	CLB_6_3_IN_pin_9_driver_mux_fanins <= track_6_3_chanY_n15 & track_6_3_chanY_n14 & track_6_3_chanY_n7 & track_6_3_chanY_n6;
	CLB_6_4_IN_pin_0_driver_mux_fanins <= track_6_4_chanX_n9 & track_6_4_chanX_n8 & track_6_4_chanX_n1 & track_6_4_chanX_n0;
	CLB_6_4_IN_pin_1_driver_mux_fanins <= track_6_4_chanY_n9 & track_6_4_chanY_n8 & track_6_4_chanY_n1 & track_6_4_chanY_n0;
	CLB_6_4_IN_pin_2_driver_mux_fanins <= track_6_3_chanX_n9 & track_6_3_chanX_n8 & track_6_3_chanX_n1 & track_6_3_chanX_n0;
	CLB_6_4_IN_pin_3_driver_mux_fanins <= track_5_4_chanY_n11 & track_5_4_chanY_n10 & track_5_4_chanY_n3 & track_5_4_chanY_n2;
	CLB_6_4_IN_pin_4_driver_mux_fanins <= track_6_4_chanX_n11 & track_6_4_chanX_n10 & track_6_4_chanX_n3 & track_6_4_chanX_n2;
	CLB_6_4_IN_pin_5_driver_mux_fanins <= track_6_4_chanY_n13 & track_6_4_chanY_n12 & track_6_4_chanY_n5 & track_6_4_chanY_n4;
	CLB_6_4_IN_pin_6_driver_mux_fanins <= track_6_3_chanX_n13 & track_6_3_chanX_n12 & track_6_3_chanX_n5 & track_6_3_chanX_n4;
	CLB_6_4_IN_pin_7_driver_mux_fanins <= track_5_4_chanY_n13 & track_5_4_chanY_n12 & track_5_4_chanY_n5 & track_5_4_chanY_n4;
	CLB_6_4_IN_pin_8_driver_mux_fanins <= track_6_4_chanX_n15 & track_6_4_chanX_n14 & track_6_4_chanX_n7 & track_6_4_chanX_n6;
	CLB_6_4_IN_pin_9_driver_mux_fanins <= track_6_4_chanY_n15 & track_6_4_chanY_n14 & track_6_4_chanY_n7 & track_6_4_chanY_n6;
	CLB_6_5_IN_pin_0_driver_mux_fanins <= track_6_5_chanX_n9 & track_6_5_chanX_n8 & track_6_5_chanX_n1 & track_6_5_chanX_n0;
	CLB_6_5_IN_pin_1_driver_mux_fanins <= track_6_5_chanY_n9 & track_6_5_chanY_n8 & track_6_5_chanY_n1 & track_6_5_chanY_n0;
	CLB_6_5_IN_pin_2_driver_mux_fanins <= track_6_4_chanX_n9 & track_6_4_chanX_n8 & track_6_4_chanX_n1 & track_6_4_chanX_n0;
	CLB_6_5_IN_pin_3_driver_mux_fanins <= track_5_5_chanY_n11 & track_5_5_chanY_n10 & track_5_5_chanY_n3 & track_5_5_chanY_n2;
	CLB_6_5_IN_pin_4_driver_mux_fanins <= track_6_5_chanX_n11 & track_6_5_chanX_n10 & track_6_5_chanX_n3 & track_6_5_chanX_n2;
	CLB_6_5_IN_pin_5_driver_mux_fanins <= track_6_5_chanY_n13 & track_6_5_chanY_n12 & track_6_5_chanY_n5 & track_6_5_chanY_n4;
	CLB_6_5_IN_pin_6_driver_mux_fanins <= track_6_4_chanX_n13 & track_6_4_chanX_n12 & track_6_4_chanX_n5 & track_6_4_chanX_n4;
	CLB_6_5_IN_pin_7_driver_mux_fanins <= track_5_5_chanY_n13 & track_5_5_chanY_n12 & track_5_5_chanY_n5 & track_5_5_chanY_n4;
	CLB_6_5_IN_pin_8_driver_mux_fanins <= track_6_5_chanX_n15 & track_6_5_chanX_n14 & track_6_5_chanX_n7 & track_6_5_chanX_n6;
	CLB_6_5_IN_pin_9_driver_mux_fanins <= track_6_5_chanY_n15 & track_6_5_chanY_n14 & track_6_5_chanY_n7 & track_6_5_chanY_n6;
	CLB_6_6_IN_pin_0_driver_mux_fanins <= track_6_6_chanX_n9 & track_6_6_chanX_n8 & track_6_6_chanX_n1 & track_6_6_chanX_n0;
	CLB_6_6_IN_pin_1_driver_mux_fanins <= track_6_6_chanY_n9 & track_6_6_chanY_n8 & track_6_6_chanY_n1 & track_6_6_chanY_n0;
	CLB_6_6_IN_pin_2_driver_mux_fanins <= track_6_5_chanX_n9 & track_6_5_chanX_n8 & track_6_5_chanX_n1 & track_6_5_chanX_n0;
	CLB_6_6_IN_pin_3_driver_mux_fanins <= track_5_6_chanY_n11 & track_5_6_chanY_n10 & track_5_6_chanY_n3 & track_5_6_chanY_n2;
	CLB_6_6_IN_pin_4_driver_mux_fanins <= track_6_6_chanX_n11 & track_6_6_chanX_n10 & track_6_6_chanX_n3 & track_6_6_chanX_n2;
	CLB_6_6_IN_pin_5_driver_mux_fanins <= track_6_6_chanY_n13 & track_6_6_chanY_n12 & track_6_6_chanY_n5 & track_6_6_chanY_n4;
	CLB_6_6_IN_pin_6_driver_mux_fanins <= track_6_5_chanX_n13 & track_6_5_chanX_n12 & track_6_5_chanX_n5 & track_6_5_chanX_n4;
	CLB_6_6_IN_pin_7_driver_mux_fanins <= track_5_6_chanY_n13 & track_5_6_chanY_n12 & track_5_6_chanY_n5 & track_5_6_chanY_n4;
	CLB_6_6_IN_pin_8_driver_mux_fanins <= track_6_6_chanX_n15 & track_6_6_chanX_n14 & track_6_6_chanX_n7 & track_6_6_chanX_n6;
	CLB_6_6_IN_pin_9_driver_mux_fanins <= track_6_6_chanY_n15 & track_6_6_chanY_n14 & track_6_6_chanY_n7 & track_6_6_chanY_n6;
	CLB_7_1_IN_pin_0_driver_mux_fanins <= track_7_1_chanX_n9 & track_7_1_chanX_n8 & track_7_1_chanX_n1 & track_7_1_chanX_n0;
	CLB_7_1_IN_pin_1_driver_mux_fanins <= track_7_1_chanY_n9 & track_7_1_chanY_n8 & track_7_1_chanY_n1 & track_7_1_chanY_n0;
	CLB_7_1_IN_pin_2_driver_mux_fanins <= track_7_0_chanX_n9 & track_7_0_chanX_n8 & track_7_0_chanX_n1 & track_7_0_chanX_n0;
	CLB_7_1_IN_pin_3_driver_mux_fanins <= track_6_1_chanY_n11 & track_6_1_chanY_n10 & track_6_1_chanY_n3 & track_6_1_chanY_n2;
	CLB_7_1_IN_pin_4_driver_mux_fanins <= track_7_1_chanX_n11 & track_7_1_chanX_n10 & track_7_1_chanX_n3 & track_7_1_chanX_n2;
	CLB_7_1_IN_pin_5_driver_mux_fanins <= track_7_1_chanY_n13 & track_7_1_chanY_n12 & track_7_1_chanY_n5 & track_7_1_chanY_n4;
	CLB_7_1_IN_pin_6_driver_mux_fanins <= track_7_0_chanX_n13 & track_7_0_chanX_n12 & track_7_0_chanX_n5 & track_7_0_chanX_n4;
	CLB_7_1_IN_pin_7_driver_mux_fanins <= track_6_1_chanY_n13 & track_6_1_chanY_n12 & track_6_1_chanY_n5 & track_6_1_chanY_n4;
	CLB_7_1_IN_pin_8_driver_mux_fanins <= track_7_1_chanX_n15 & track_7_1_chanX_n14 & track_7_1_chanX_n7 & track_7_1_chanX_n6;
	CLB_7_1_IN_pin_9_driver_mux_fanins <= track_7_1_chanY_n15 & track_7_1_chanY_n14 & track_7_1_chanY_n7 & track_7_1_chanY_n6;
	CLB_7_2_IN_pin_0_driver_mux_fanins <= track_7_2_chanX_n9 & track_7_2_chanX_n8 & track_7_2_chanX_n1 & track_7_2_chanX_n0;
	CLB_7_2_IN_pin_1_driver_mux_fanins <= track_7_2_chanY_n9 & track_7_2_chanY_n8 & track_7_2_chanY_n1 & track_7_2_chanY_n0;
	CLB_7_2_IN_pin_2_driver_mux_fanins <= track_7_1_chanX_n9 & track_7_1_chanX_n8 & track_7_1_chanX_n1 & track_7_1_chanX_n0;
	CLB_7_2_IN_pin_3_driver_mux_fanins <= track_6_2_chanY_n11 & track_6_2_chanY_n10 & track_6_2_chanY_n3 & track_6_2_chanY_n2;
	CLB_7_2_IN_pin_4_driver_mux_fanins <= track_7_2_chanX_n11 & track_7_2_chanX_n10 & track_7_2_chanX_n3 & track_7_2_chanX_n2;
	CLB_7_2_IN_pin_5_driver_mux_fanins <= track_7_2_chanY_n13 & track_7_2_chanY_n12 & track_7_2_chanY_n5 & track_7_2_chanY_n4;
	CLB_7_2_IN_pin_6_driver_mux_fanins <= track_7_1_chanX_n13 & track_7_1_chanX_n12 & track_7_1_chanX_n5 & track_7_1_chanX_n4;
	CLB_7_2_IN_pin_7_driver_mux_fanins <= track_6_2_chanY_n13 & track_6_2_chanY_n12 & track_6_2_chanY_n5 & track_6_2_chanY_n4;
	CLB_7_2_IN_pin_8_driver_mux_fanins <= track_7_2_chanX_n15 & track_7_2_chanX_n14 & track_7_2_chanX_n7 & track_7_2_chanX_n6;
	CLB_7_2_IN_pin_9_driver_mux_fanins <= track_7_2_chanY_n15 & track_7_2_chanY_n14 & track_7_2_chanY_n7 & track_7_2_chanY_n6;
	CLB_7_3_IN_pin_0_driver_mux_fanins <= track_7_3_chanX_n9 & track_7_3_chanX_n8 & track_7_3_chanX_n1 & track_7_3_chanX_n0;
	CLB_7_3_IN_pin_1_driver_mux_fanins <= track_7_3_chanY_n9 & track_7_3_chanY_n8 & track_7_3_chanY_n1 & track_7_3_chanY_n0;
	CLB_7_3_IN_pin_2_driver_mux_fanins <= track_7_2_chanX_n9 & track_7_2_chanX_n8 & track_7_2_chanX_n1 & track_7_2_chanX_n0;
	CLB_7_3_IN_pin_3_driver_mux_fanins <= track_6_3_chanY_n11 & track_6_3_chanY_n10 & track_6_3_chanY_n3 & track_6_3_chanY_n2;
	CLB_7_3_IN_pin_4_driver_mux_fanins <= track_7_3_chanX_n11 & track_7_3_chanX_n10 & track_7_3_chanX_n3 & track_7_3_chanX_n2;
	CLB_7_3_IN_pin_5_driver_mux_fanins <= track_7_3_chanY_n13 & track_7_3_chanY_n12 & track_7_3_chanY_n5 & track_7_3_chanY_n4;
	CLB_7_3_IN_pin_6_driver_mux_fanins <= track_7_2_chanX_n13 & track_7_2_chanX_n12 & track_7_2_chanX_n5 & track_7_2_chanX_n4;
	CLB_7_3_IN_pin_7_driver_mux_fanins <= track_6_3_chanY_n13 & track_6_3_chanY_n12 & track_6_3_chanY_n5 & track_6_3_chanY_n4;
	CLB_7_3_IN_pin_8_driver_mux_fanins <= track_7_3_chanX_n15 & track_7_3_chanX_n14 & track_7_3_chanX_n7 & track_7_3_chanX_n6;
	CLB_7_3_IN_pin_9_driver_mux_fanins <= track_7_3_chanY_n15 & track_7_3_chanY_n14 & track_7_3_chanY_n7 & track_7_3_chanY_n6;
	CLB_7_4_IN_pin_0_driver_mux_fanins <= track_7_4_chanX_n9 & track_7_4_chanX_n8 & track_7_4_chanX_n1 & track_7_4_chanX_n0;
	CLB_7_4_IN_pin_1_driver_mux_fanins <= track_7_4_chanY_n9 & track_7_4_chanY_n8 & track_7_4_chanY_n1 & track_7_4_chanY_n0;
	CLB_7_4_IN_pin_2_driver_mux_fanins <= track_7_3_chanX_n9 & track_7_3_chanX_n8 & track_7_3_chanX_n1 & track_7_3_chanX_n0;
	CLB_7_4_IN_pin_3_driver_mux_fanins <= track_6_4_chanY_n11 & track_6_4_chanY_n10 & track_6_4_chanY_n3 & track_6_4_chanY_n2;
	CLB_7_4_IN_pin_4_driver_mux_fanins <= track_7_4_chanX_n11 & track_7_4_chanX_n10 & track_7_4_chanX_n3 & track_7_4_chanX_n2;
	CLB_7_4_IN_pin_5_driver_mux_fanins <= track_7_4_chanY_n13 & track_7_4_chanY_n12 & track_7_4_chanY_n5 & track_7_4_chanY_n4;
	CLB_7_4_IN_pin_6_driver_mux_fanins <= track_7_3_chanX_n13 & track_7_3_chanX_n12 & track_7_3_chanX_n5 & track_7_3_chanX_n4;
	CLB_7_4_IN_pin_7_driver_mux_fanins <= track_6_4_chanY_n13 & track_6_4_chanY_n12 & track_6_4_chanY_n5 & track_6_4_chanY_n4;
	CLB_7_4_IN_pin_8_driver_mux_fanins <= track_7_4_chanX_n15 & track_7_4_chanX_n14 & track_7_4_chanX_n7 & track_7_4_chanX_n6;
	CLB_7_4_IN_pin_9_driver_mux_fanins <= track_7_4_chanY_n15 & track_7_4_chanY_n14 & track_7_4_chanY_n7 & track_7_4_chanY_n6;
	CLB_7_5_IN_pin_0_driver_mux_fanins <= track_7_5_chanX_n9 & track_7_5_chanX_n8 & track_7_5_chanX_n1 & track_7_5_chanX_n0;
	CLB_7_5_IN_pin_1_driver_mux_fanins <= track_7_5_chanY_n9 & track_7_5_chanY_n8 & track_7_5_chanY_n1 & track_7_5_chanY_n0;
	CLB_7_5_IN_pin_2_driver_mux_fanins <= track_7_4_chanX_n9 & track_7_4_chanX_n8 & track_7_4_chanX_n1 & track_7_4_chanX_n0;
	CLB_7_5_IN_pin_3_driver_mux_fanins <= track_6_5_chanY_n11 & track_6_5_chanY_n10 & track_6_5_chanY_n3 & track_6_5_chanY_n2;
	CLB_7_5_IN_pin_4_driver_mux_fanins <= track_7_5_chanX_n11 & track_7_5_chanX_n10 & track_7_5_chanX_n3 & track_7_5_chanX_n2;
	CLB_7_5_IN_pin_5_driver_mux_fanins <= track_7_5_chanY_n13 & track_7_5_chanY_n12 & track_7_5_chanY_n5 & track_7_5_chanY_n4;
	CLB_7_5_IN_pin_6_driver_mux_fanins <= track_7_4_chanX_n13 & track_7_4_chanX_n12 & track_7_4_chanX_n5 & track_7_4_chanX_n4;
	CLB_7_5_IN_pin_7_driver_mux_fanins <= track_6_5_chanY_n13 & track_6_5_chanY_n12 & track_6_5_chanY_n5 & track_6_5_chanY_n4;
	CLB_7_5_IN_pin_8_driver_mux_fanins <= track_7_5_chanX_n15 & track_7_5_chanX_n14 & track_7_5_chanX_n7 & track_7_5_chanX_n6;
	CLB_7_5_IN_pin_9_driver_mux_fanins <= track_7_5_chanY_n15 & track_7_5_chanY_n14 & track_7_5_chanY_n7 & track_7_5_chanY_n6;
	CLB_7_6_IN_pin_0_driver_mux_fanins <= track_7_6_chanX_n9 & track_7_6_chanX_n8 & track_7_6_chanX_n1 & track_7_6_chanX_n0;
	CLB_7_6_IN_pin_1_driver_mux_fanins <= track_7_6_chanY_n9 & track_7_6_chanY_n8 & track_7_6_chanY_n1 & track_7_6_chanY_n0;
	CLB_7_6_IN_pin_2_driver_mux_fanins <= track_7_5_chanX_n9 & track_7_5_chanX_n8 & track_7_5_chanX_n1 & track_7_5_chanX_n0;
	CLB_7_6_IN_pin_3_driver_mux_fanins <= track_6_6_chanY_n11 & track_6_6_chanY_n10 & track_6_6_chanY_n3 & track_6_6_chanY_n2;
	CLB_7_6_IN_pin_4_driver_mux_fanins <= track_7_6_chanX_n11 & track_7_6_chanX_n10 & track_7_6_chanX_n3 & track_7_6_chanX_n2;
	CLB_7_6_IN_pin_5_driver_mux_fanins <= track_7_6_chanY_n13 & track_7_6_chanY_n12 & track_7_6_chanY_n5 & track_7_6_chanY_n4;
	CLB_7_6_IN_pin_6_driver_mux_fanins <= track_7_5_chanX_n13 & track_7_5_chanX_n12 & track_7_5_chanX_n5 & track_7_5_chanX_n4;
	CLB_7_6_IN_pin_7_driver_mux_fanins <= track_6_6_chanY_n13 & track_6_6_chanY_n12 & track_6_6_chanY_n5 & track_6_6_chanY_n4;
	CLB_7_6_IN_pin_8_driver_mux_fanins <= track_7_6_chanX_n15 & track_7_6_chanX_n14 & track_7_6_chanX_n7 & track_7_6_chanX_n6;
	CLB_7_6_IN_pin_9_driver_mux_fanins <= track_7_6_chanY_n15 & track_7_6_chanY_n14 & track_7_6_chanY_n7 & track_7_6_chanY_n6;
	CLB_8_1_IN_pin_0_driver_mux_fanins <= track_8_1_chanX_n9 & track_8_1_chanX_n8 & track_8_1_chanX_n1 & track_8_1_chanX_n0;
	CLB_8_1_IN_pin_1_driver_mux_fanins <= track_8_1_chanY_n9 & track_8_1_chanY_n8 & track_8_1_chanY_n1 & track_8_1_chanY_n0;
	CLB_8_1_IN_pin_2_driver_mux_fanins <= track_8_0_chanX_n9 & track_8_0_chanX_n8 & track_8_0_chanX_n1 & track_8_0_chanX_n0;
	CLB_8_1_IN_pin_3_driver_mux_fanins <= track_7_1_chanY_n11 & track_7_1_chanY_n10 & track_7_1_chanY_n3 & track_7_1_chanY_n2;
	CLB_8_1_IN_pin_4_driver_mux_fanins <= track_8_1_chanX_n11 & track_8_1_chanX_n10 & track_8_1_chanX_n3 & track_8_1_chanX_n2;
	CLB_8_1_IN_pin_5_driver_mux_fanins <= track_8_1_chanY_n13 & track_8_1_chanY_n12 & track_8_1_chanY_n5 & track_8_1_chanY_n4;
	CLB_8_1_IN_pin_6_driver_mux_fanins <= track_8_0_chanX_n13 & track_8_0_chanX_n12 & track_8_0_chanX_n5 & track_8_0_chanX_n4;
	CLB_8_1_IN_pin_7_driver_mux_fanins <= track_7_1_chanY_n13 & track_7_1_chanY_n12 & track_7_1_chanY_n5 & track_7_1_chanY_n4;
	CLB_8_1_IN_pin_8_driver_mux_fanins <= track_8_1_chanX_n15 & track_8_1_chanX_n14 & track_8_1_chanX_n7 & track_8_1_chanX_n6;
	CLB_8_1_IN_pin_9_driver_mux_fanins <= track_8_1_chanY_n15 & track_8_1_chanY_n14 & track_8_1_chanY_n7 & track_8_1_chanY_n6;
	CLB_8_2_IN_pin_0_driver_mux_fanins <= track_8_2_chanX_n9 & track_8_2_chanX_n8 & track_8_2_chanX_n1 & track_8_2_chanX_n0;
	CLB_8_2_IN_pin_1_driver_mux_fanins <= track_8_2_chanY_n9 & track_8_2_chanY_n8 & track_8_2_chanY_n1 & track_8_2_chanY_n0;
	CLB_8_2_IN_pin_2_driver_mux_fanins <= track_8_1_chanX_n9 & track_8_1_chanX_n8 & track_8_1_chanX_n1 & track_8_1_chanX_n0;
	CLB_8_2_IN_pin_3_driver_mux_fanins <= track_7_2_chanY_n11 & track_7_2_chanY_n10 & track_7_2_chanY_n3 & track_7_2_chanY_n2;
	CLB_8_2_IN_pin_4_driver_mux_fanins <= track_8_2_chanX_n11 & track_8_2_chanX_n10 & track_8_2_chanX_n3 & track_8_2_chanX_n2;
	CLB_8_2_IN_pin_5_driver_mux_fanins <= track_8_2_chanY_n13 & track_8_2_chanY_n12 & track_8_2_chanY_n5 & track_8_2_chanY_n4;
	CLB_8_2_IN_pin_6_driver_mux_fanins <= track_8_1_chanX_n13 & track_8_1_chanX_n12 & track_8_1_chanX_n5 & track_8_1_chanX_n4;
	CLB_8_2_IN_pin_7_driver_mux_fanins <= track_7_2_chanY_n13 & track_7_2_chanY_n12 & track_7_2_chanY_n5 & track_7_2_chanY_n4;
	CLB_8_2_IN_pin_8_driver_mux_fanins <= track_8_2_chanX_n15 & track_8_2_chanX_n14 & track_8_2_chanX_n7 & track_8_2_chanX_n6;
	CLB_8_2_IN_pin_9_driver_mux_fanins <= track_8_2_chanY_n15 & track_8_2_chanY_n14 & track_8_2_chanY_n7 & track_8_2_chanY_n6;
	CLB_8_3_IN_pin_0_driver_mux_fanins <= track_8_3_chanX_n9 & track_8_3_chanX_n8 & track_8_3_chanX_n1 & track_8_3_chanX_n0;
	CLB_8_3_IN_pin_1_driver_mux_fanins <= track_8_3_chanY_n9 & track_8_3_chanY_n8 & track_8_3_chanY_n1 & track_8_3_chanY_n0;
	CLB_8_3_IN_pin_2_driver_mux_fanins <= track_8_2_chanX_n9 & track_8_2_chanX_n8 & track_8_2_chanX_n1 & track_8_2_chanX_n0;
	CLB_8_3_IN_pin_3_driver_mux_fanins <= track_7_3_chanY_n11 & track_7_3_chanY_n10 & track_7_3_chanY_n3 & track_7_3_chanY_n2;
	CLB_8_3_IN_pin_4_driver_mux_fanins <= track_8_3_chanX_n11 & track_8_3_chanX_n10 & track_8_3_chanX_n3 & track_8_3_chanX_n2;
	CLB_8_3_IN_pin_5_driver_mux_fanins <= track_8_3_chanY_n13 & track_8_3_chanY_n12 & track_8_3_chanY_n5 & track_8_3_chanY_n4;
	CLB_8_3_IN_pin_6_driver_mux_fanins <= track_8_2_chanX_n13 & track_8_2_chanX_n12 & track_8_2_chanX_n5 & track_8_2_chanX_n4;
	CLB_8_3_IN_pin_7_driver_mux_fanins <= track_7_3_chanY_n13 & track_7_3_chanY_n12 & track_7_3_chanY_n5 & track_7_3_chanY_n4;
	CLB_8_3_IN_pin_8_driver_mux_fanins <= track_8_3_chanX_n15 & track_8_3_chanX_n14 & track_8_3_chanX_n7 & track_8_3_chanX_n6;
	CLB_8_3_IN_pin_9_driver_mux_fanins <= track_8_3_chanY_n15 & track_8_3_chanY_n14 & track_8_3_chanY_n7 & track_8_3_chanY_n6;
	CLB_8_4_IN_pin_0_driver_mux_fanins <= track_8_4_chanX_n9 & track_8_4_chanX_n8 & track_8_4_chanX_n1 & track_8_4_chanX_n0;
	CLB_8_4_IN_pin_1_driver_mux_fanins <= track_8_4_chanY_n9 & track_8_4_chanY_n8 & track_8_4_chanY_n1 & track_8_4_chanY_n0;
	CLB_8_4_IN_pin_2_driver_mux_fanins <= track_8_3_chanX_n9 & track_8_3_chanX_n8 & track_8_3_chanX_n1 & track_8_3_chanX_n0;
	CLB_8_4_IN_pin_3_driver_mux_fanins <= track_7_4_chanY_n11 & track_7_4_chanY_n10 & track_7_4_chanY_n3 & track_7_4_chanY_n2;
	CLB_8_4_IN_pin_4_driver_mux_fanins <= track_8_4_chanX_n11 & track_8_4_chanX_n10 & track_8_4_chanX_n3 & track_8_4_chanX_n2;
	CLB_8_4_IN_pin_5_driver_mux_fanins <= track_8_4_chanY_n13 & track_8_4_chanY_n12 & track_8_4_chanY_n5 & track_8_4_chanY_n4;
	CLB_8_4_IN_pin_6_driver_mux_fanins <= track_8_3_chanX_n13 & track_8_3_chanX_n12 & track_8_3_chanX_n5 & track_8_3_chanX_n4;
	CLB_8_4_IN_pin_7_driver_mux_fanins <= track_7_4_chanY_n13 & track_7_4_chanY_n12 & track_7_4_chanY_n5 & track_7_4_chanY_n4;
	CLB_8_4_IN_pin_8_driver_mux_fanins <= track_8_4_chanX_n15 & track_8_4_chanX_n14 & track_8_4_chanX_n7 & track_8_4_chanX_n6;
	CLB_8_4_IN_pin_9_driver_mux_fanins <= track_8_4_chanY_n15 & track_8_4_chanY_n14 & track_8_4_chanY_n7 & track_8_4_chanY_n6;
	CLB_8_5_IN_pin_0_driver_mux_fanins <= track_8_5_chanX_n9 & track_8_5_chanX_n8 & track_8_5_chanX_n1 & track_8_5_chanX_n0;
	CLB_8_5_IN_pin_1_driver_mux_fanins <= track_8_5_chanY_n9 & track_8_5_chanY_n8 & track_8_5_chanY_n1 & track_8_5_chanY_n0;
	CLB_8_5_IN_pin_2_driver_mux_fanins <= track_8_4_chanX_n9 & track_8_4_chanX_n8 & track_8_4_chanX_n1 & track_8_4_chanX_n0;
	CLB_8_5_IN_pin_3_driver_mux_fanins <= track_7_5_chanY_n11 & track_7_5_chanY_n10 & track_7_5_chanY_n3 & track_7_5_chanY_n2;
	CLB_8_5_IN_pin_4_driver_mux_fanins <= track_8_5_chanX_n11 & track_8_5_chanX_n10 & track_8_5_chanX_n3 & track_8_5_chanX_n2;
	CLB_8_5_IN_pin_5_driver_mux_fanins <= track_8_5_chanY_n13 & track_8_5_chanY_n12 & track_8_5_chanY_n5 & track_8_5_chanY_n4;
	CLB_8_5_IN_pin_6_driver_mux_fanins <= track_8_4_chanX_n13 & track_8_4_chanX_n12 & track_8_4_chanX_n5 & track_8_4_chanX_n4;
	CLB_8_5_IN_pin_7_driver_mux_fanins <= track_7_5_chanY_n13 & track_7_5_chanY_n12 & track_7_5_chanY_n5 & track_7_5_chanY_n4;
	CLB_8_5_IN_pin_8_driver_mux_fanins <= track_8_5_chanX_n15 & track_8_5_chanX_n14 & track_8_5_chanX_n7 & track_8_5_chanX_n6;
	CLB_8_5_IN_pin_9_driver_mux_fanins <= track_8_5_chanY_n15 & track_8_5_chanY_n14 & track_8_5_chanY_n7 & track_8_5_chanY_n6;
	CLB_8_6_IN_pin_0_driver_mux_fanins <= track_8_6_chanX_n9 & track_8_6_chanX_n8 & track_8_6_chanX_n1 & track_8_6_chanX_n0;
	CLB_8_6_IN_pin_1_driver_mux_fanins <= track_8_6_chanY_n9 & track_8_6_chanY_n8 & track_8_6_chanY_n1 & track_8_6_chanY_n0;
	CLB_8_6_IN_pin_2_driver_mux_fanins <= track_8_5_chanX_n9 & track_8_5_chanX_n8 & track_8_5_chanX_n1 & track_8_5_chanX_n0;
	CLB_8_6_IN_pin_3_driver_mux_fanins <= track_7_6_chanY_n11 & track_7_6_chanY_n10 & track_7_6_chanY_n3 & track_7_6_chanY_n2;
	CLB_8_6_IN_pin_4_driver_mux_fanins <= track_8_6_chanX_n11 & track_8_6_chanX_n10 & track_8_6_chanX_n3 & track_8_6_chanX_n2;
	CLB_8_6_IN_pin_5_driver_mux_fanins <= track_8_6_chanY_n13 & track_8_6_chanY_n12 & track_8_6_chanY_n5 & track_8_6_chanY_n4;
	CLB_8_6_IN_pin_6_driver_mux_fanins <= track_8_5_chanX_n13 & track_8_5_chanX_n12 & track_8_5_chanX_n5 & track_8_5_chanX_n4;
	CLB_8_6_IN_pin_7_driver_mux_fanins <= track_7_6_chanY_n13 & track_7_6_chanY_n12 & track_7_6_chanY_n5 & track_7_6_chanY_n4;
	CLB_8_6_IN_pin_8_driver_mux_fanins <= track_8_6_chanX_n15 & track_8_6_chanX_n14 & track_8_6_chanX_n7 & track_8_6_chanX_n6;
	CLB_8_6_IN_pin_9_driver_mux_fanins <= track_8_6_chanY_n15 & track_8_6_chanY_n14 & track_8_6_chanY_n7 & track_8_6_chanY_n6;
	IO_0_1_IN_pin_0_driver_mux_fanins  <= track_0_1_chanY_n13 & track_0_1_chanY_n12 & track_0_1_chanY_n9 & track_0_1_chanY_n8 & track_0_1_chanY_n5 & track_0_1_chanY_n4 & track_0_1_chanY_n1 & track_0_1_chanY_n0;
	IO_0_1_IN_pin_1_driver_mux_fanins  <= track_0_1_chanY_n15 & track_0_1_chanY_n14 & track_0_1_chanY_n11 & track_0_1_chanY_n10 & track_0_1_chanY_n7 & track_0_1_chanY_n6 & track_0_1_chanY_n3 & track_0_1_chanY_n2;
	IO_0_2_IN_pin_0_driver_mux_fanins  <= track_0_2_chanY_n13 & track_0_2_chanY_n12 & track_0_2_chanY_n9 & track_0_2_chanY_n8 & track_0_2_chanY_n5 & track_0_2_chanY_n4 & track_0_2_chanY_n1 & track_0_2_chanY_n0;
	IO_0_2_IN_pin_1_driver_mux_fanins  <= track_0_2_chanY_n15 & track_0_2_chanY_n14 & track_0_2_chanY_n11 & track_0_2_chanY_n10 & track_0_2_chanY_n7 & track_0_2_chanY_n6 & track_0_2_chanY_n3 & track_0_2_chanY_n2;
	IO_0_3_IN_pin_0_driver_mux_fanins  <= track_0_3_chanY_n13 & track_0_3_chanY_n12 & track_0_3_chanY_n9 & track_0_3_chanY_n8 & track_0_3_chanY_n5 & track_0_3_chanY_n4 & track_0_3_chanY_n1 & track_0_3_chanY_n0;
	IO_0_3_IN_pin_1_driver_mux_fanins  <= track_0_3_chanY_n15 & track_0_3_chanY_n14 & track_0_3_chanY_n11 & track_0_3_chanY_n10 & track_0_3_chanY_n7 & track_0_3_chanY_n6 & track_0_3_chanY_n3 & track_0_3_chanY_n2;
	IO_0_4_IN_pin_0_driver_mux_fanins  <= track_0_4_chanY_n13 & track_0_4_chanY_n12 & track_0_4_chanY_n9 & track_0_4_chanY_n8 & track_0_4_chanY_n5 & track_0_4_chanY_n4 & track_0_4_chanY_n1 & track_0_4_chanY_n0;
	IO_0_4_IN_pin_1_driver_mux_fanins  <= track_0_4_chanY_n15 & track_0_4_chanY_n14 & track_0_4_chanY_n11 & track_0_4_chanY_n10 & track_0_4_chanY_n7 & track_0_4_chanY_n6 & track_0_4_chanY_n3 & track_0_4_chanY_n2;
	IO_0_5_IN_pin_0_driver_mux_fanins  <= track_0_5_chanY_n13 & track_0_5_chanY_n12 & track_0_5_chanY_n9 & track_0_5_chanY_n8 & track_0_5_chanY_n5 & track_0_5_chanY_n4 & track_0_5_chanY_n1 & track_0_5_chanY_n0;
	IO_0_5_IN_pin_1_driver_mux_fanins  <= track_0_5_chanY_n15 & track_0_5_chanY_n14 & track_0_5_chanY_n11 & track_0_5_chanY_n10 & track_0_5_chanY_n7 & track_0_5_chanY_n6 & track_0_5_chanY_n3 & track_0_5_chanY_n2;
	IO_0_6_IN_pin_0_driver_mux_fanins  <= track_0_6_chanY_n13 & track_0_6_chanY_n12 & track_0_6_chanY_n9 & track_0_6_chanY_n8 & track_0_6_chanY_n5 & track_0_6_chanY_n4 & track_0_6_chanY_n1 & track_0_6_chanY_n0;
	IO_0_6_IN_pin_1_driver_mux_fanins  <= track_0_6_chanY_n15 & track_0_6_chanY_n14 & track_0_6_chanY_n11 & track_0_6_chanY_n10 & track_0_6_chanY_n7 & track_0_6_chanY_n6 & track_0_6_chanY_n3 & track_0_6_chanY_n2;
	IO_1_0_IN_pin_0_driver_mux_fanins  <= track_1_0_chanX_n13 & track_1_0_chanX_n12 & track_1_0_chanX_n9 & track_1_0_chanX_n8 & track_1_0_chanX_n5 & track_1_0_chanX_n4 & track_1_0_chanX_n1 & track_1_0_chanX_n0;
	IO_1_0_IN_pin_1_driver_mux_fanins  <= track_1_0_chanX_n15 & track_1_0_chanX_n14 & track_1_0_chanX_n11 & track_1_0_chanX_n10 & track_1_0_chanX_n7 & track_1_0_chanX_n6 & track_1_0_chanX_n3 & track_1_0_chanX_n2;
	IO_1_7_IN_pin_0_driver_mux_fanins  <= track_1_6_chanX_n13 & track_1_6_chanX_n12 & track_1_6_chanX_n9 & track_1_6_chanX_n8 & track_1_6_chanX_n5 & track_1_6_chanX_n4 & track_1_6_chanX_n1 & track_1_6_chanX_n0;
	IO_1_7_IN_pin_1_driver_mux_fanins  <= track_1_6_chanX_n15 & track_1_6_chanX_n14 & track_1_6_chanX_n11 & track_1_6_chanX_n10 & track_1_6_chanX_n7 & track_1_6_chanX_n6 & track_1_6_chanX_n3 & track_1_6_chanX_n2;
	IO_2_0_IN_pin_0_driver_mux_fanins  <= track_2_0_chanX_n13 & track_2_0_chanX_n12 & track_2_0_chanX_n9 & track_2_0_chanX_n8 & track_2_0_chanX_n5 & track_2_0_chanX_n4 & track_2_0_chanX_n1 & track_2_0_chanX_n0;
	IO_2_0_IN_pin_1_driver_mux_fanins  <= track_2_0_chanX_n15 & track_2_0_chanX_n14 & track_2_0_chanX_n11 & track_2_0_chanX_n10 & track_2_0_chanX_n7 & track_2_0_chanX_n6 & track_2_0_chanX_n3 & track_2_0_chanX_n2;
	IO_2_7_IN_pin_0_driver_mux_fanins  <= track_2_6_chanX_n13 & track_2_6_chanX_n12 & track_2_6_chanX_n9 & track_2_6_chanX_n8 & track_2_6_chanX_n5 & track_2_6_chanX_n4 & track_2_6_chanX_n1 & track_2_6_chanX_n0;
	IO_2_7_IN_pin_1_driver_mux_fanins  <= track_2_6_chanX_n15 & track_2_6_chanX_n14 & track_2_6_chanX_n11 & track_2_6_chanX_n10 & track_2_6_chanX_n7 & track_2_6_chanX_n6 & track_2_6_chanX_n3 & track_2_6_chanX_n2;
	IO_3_0_IN_pin_0_driver_mux_fanins  <= track_3_0_chanX_n13 & track_3_0_chanX_n12 & track_3_0_chanX_n9 & track_3_0_chanX_n8 & track_3_0_chanX_n5 & track_3_0_chanX_n4 & track_3_0_chanX_n1 & track_3_0_chanX_n0;
	IO_3_0_IN_pin_1_driver_mux_fanins  <= track_3_0_chanX_n15 & track_3_0_chanX_n14 & track_3_0_chanX_n11 & track_3_0_chanX_n10 & track_3_0_chanX_n7 & track_3_0_chanX_n6 & track_3_0_chanX_n3 & track_3_0_chanX_n2;
	IO_3_7_IN_pin_0_driver_mux_fanins  <= track_3_6_chanX_n13 & track_3_6_chanX_n12 & track_3_6_chanX_n9 & track_3_6_chanX_n8 & track_3_6_chanX_n5 & track_3_6_chanX_n4 & track_3_6_chanX_n1 & track_3_6_chanX_n0;
	IO_3_7_IN_pin_1_driver_mux_fanins  <= track_3_6_chanX_n15 & track_3_6_chanX_n14 & track_3_6_chanX_n11 & track_3_6_chanX_n10 & track_3_6_chanX_n7 & track_3_6_chanX_n6 & track_3_6_chanX_n3 & track_3_6_chanX_n2;
	IO_4_0_IN_pin_0_driver_mux_fanins  <= track_4_0_chanX_n13 & track_4_0_chanX_n12 & track_4_0_chanX_n9 & track_4_0_chanX_n8 & track_4_0_chanX_n5 & track_4_0_chanX_n4 & track_4_0_chanX_n1 & track_4_0_chanX_n0;
	IO_4_0_IN_pin_1_driver_mux_fanins  <= track_4_0_chanX_n15 & track_4_0_chanX_n14 & track_4_0_chanX_n11 & track_4_0_chanX_n10 & track_4_0_chanX_n7 & track_4_0_chanX_n6 & track_4_0_chanX_n3 & track_4_0_chanX_n2;
	IO_4_7_IN_pin_0_driver_mux_fanins  <= track_4_6_chanX_n13 & track_4_6_chanX_n12 & track_4_6_chanX_n9 & track_4_6_chanX_n8 & track_4_6_chanX_n5 & track_4_6_chanX_n4 & track_4_6_chanX_n1 & track_4_6_chanX_n0;
	IO_4_7_IN_pin_1_driver_mux_fanins  <= track_4_6_chanX_n15 & track_4_6_chanX_n14 & track_4_6_chanX_n11 & track_4_6_chanX_n10 & track_4_6_chanX_n7 & track_4_6_chanX_n6 & track_4_6_chanX_n3 & track_4_6_chanX_n2;
	IO_5_0_IN_pin_0_driver_mux_fanins  <= track_5_0_chanX_n13 & track_5_0_chanX_n12 & track_5_0_chanX_n9 & track_5_0_chanX_n8 & track_5_0_chanX_n5 & track_5_0_chanX_n4 & track_5_0_chanX_n1 & track_5_0_chanX_n0;
	IO_5_0_IN_pin_1_driver_mux_fanins  <= track_5_0_chanX_n15 & track_5_0_chanX_n14 & track_5_0_chanX_n11 & track_5_0_chanX_n10 & track_5_0_chanX_n7 & track_5_0_chanX_n6 & track_5_0_chanX_n3 & track_5_0_chanX_n2;
	IO_5_7_IN_pin_0_driver_mux_fanins  <= track_5_6_chanX_n13 & track_5_6_chanX_n12 & track_5_6_chanX_n9 & track_5_6_chanX_n8 & track_5_6_chanX_n5 & track_5_6_chanX_n4 & track_5_6_chanX_n1 & track_5_6_chanX_n0;
	IO_5_7_IN_pin_1_driver_mux_fanins  <= track_5_6_chanX_n15 & track_5_6_chanX_n14 & track_5_6_chanX_n11 & track_5_6_chanX_n10 & track_5_6_chanX_n7 & track_5_6_chanX_n6 & track_5_6_chanX_n3 & track_5_6_chanX_n2;
	IO_6_0_IN_pin_0_driver_mux_fanins  <= track_6_0_chanX_n13 & track_6_0_chanX_n12 & track_6_0_chanX_n9 & track_6_0_chanX_n8 & track_6_0_chanX_n5 & track_6_0_chanX_n4 & track_6_0_chanX_n1 & track_6_0_chanX_n0;
	IO_6_0_IN_pin_1_driver_mux_fanins  <= track_6_0_chanX_n15 & track_6_0_chanX_n14 & track_6_0_chanX_n11 & track_6_0_chanX_n10 & track_6_0_chanX_n7 & track_6_0_chanX_n6 & track_6_0_chanX_n3 & track_6_0_chanX_n2;
	IO_6_7_IN_pin_0_driver_mux_fanins  <= track_6_6_chanX_n13 & track_6_6_chanX_n12 & track_6_6_chanX_n9 & track_6_6_chanX_n8 & track_6_6_chanX_n5 & track_6_6_chanX_n4 & track_6_6_chanX_n1 & track_6_6_chanX_n0;
	IO_6_7_IN_pin_1_driver_mux_fanins  <= track_6_6_chanX_n15 & track_6_6_chanX_n14 & track_6_6_chanX_n11 & track_6_6_chanX_n10 & track_6_6_chanX_n7 & track_6_6_chanX_n6 & track_6_6_chanX_n3 & track_6_6_chanX_n2;
	IO_7_0_IN_pin_0_driver_mux_fanins  <= track_7_0_chanX_n13 & track_7_0_chanX_n12 & track_7_0_chanX_n9 & track_7_0_chanX_n8 & track_7_0_chanX_n5 & track_7_0_chanX_n4 & track_7_0_chanX_n1 & track_7_0_chanX_n0;
	IO_7_0_IN_pin_1_driver_mux_fanins  <= track_7_0_chanX_n15 & track_7_0_chanX_n14 & track_7_0_chanX_n11 & track_7_0_chanX_n10 & track_7_0_chanX_n7 & track_7_0_chanX_n6 & track_7_0_chanX_n3 & track_7_0_chanX_n2;
	IO_7_7_IN_pin_0_driver_mux_fanins  <= track_7_6_chanX_n13 & track_7_6_chanX_n12 & track_7_6_chanX_n9 & track_7_6_chanX_n8 & track_7_6_chanX_n5 & track_7_6_chanX_n4 & track_7_6_chanX_n1 & track_7_6_chanX_n0;
	IO_7_7_IN_pin_1_driver_mux_fanins  <= track_7_6_chanX_n15 & track_7_6_chanX_n14 & track_7_6_chanX_n11 & track_7_6_chanX_n10 & track_7_6_chanX_n7 & track_7_6_chanX_n6 & track_7_6_chanX_n3 & track_7_6_chanX_n2;
	IO_8_0_IN_pin_0_driver_mux_fanins  <= track_8_0_chanX_n13 & track_8_0_chanX_n12 & track_8_0_chanX_n9 & track_8_0_chanX_n8 & track_8_0_chanX_n5 & track_8_0_chanX_n4 & track_8_0_chanX_n1 & track_8_0_chanX_n0;
	IO_8_0_IN_pin_1_driver_mux_fanins  <= track_8_0_chanX_n15 & track_8_0_chanX_n14 & track_8_0_chanX_n11 & track_8_0_chanX_n10 & track_8_0_chanX_n7 & track_8_0_chanX_n6 & track_8_0_chanX_n3 & track_8_0_chanX_n2;
	IO_8_7_IN_pin_0_driver_mux_fanins  <= track_8_6_chanX_n13 & track_8_6_chanX_n12 & track_8_6_chanX_n9 & track_8_6_chanX_n8 & track_8_6_chanX_n5 & track_8_6_chanX_n4 & track_8_6_chanX_n1 & track_8_6_chanX_n0;
	IO_8_7_IN_pin_1_driver_mux_fanins  <= track_8_6_chanX_n15 & track_8_6_chanX_n14 & track_8_6_chanX_n11 & track_8_6_chanX_n10 & track_8_6_chanX_n7 & track_8_6_chanX_n6 & track_8_6_chanX_n3 & track_8_6_chanX_n2;
	IO_9_1_IN_pin_0_driver_mux_fanins  <= track_8_1_chanY_n13 & track_8_1_chanY_n12 & track_8_1_chanY_n9 & track_8_1_chanY_n8 & track_8_1_chanY_n5 & track_8_1_chanY_n4 & track_8_1_chanY_n1 & track_8_1_chanY_n0;
	IO_9_1_IN_pin_1_driver_mux_fanins  <= track_8_1_chanY_n15 & track_8_1_chanY_n14 & track_8_1_chanY_n11 & track_8_1_chanY_n10 & track_8_1_chanY_n7 & track_8_1_chanY_n6 & track_8_1_chanY_n3 & track_8_1_chanY_n2;
	IO_9_2_IN_pin_0_driver_mux_fanins  <= track_8_2_chanY_n13 & track_8_2_chanY_n12 & track_8_2_chanY_n9 & track_8_2_chanY_n8 & track_8_2_chanY_n5 & track_8_2_chanY_n4 & track_8_2_chanY_n1 & track_8_2_chanY_n0;
	IO_9_2_IN_pin_1_driver_mux_fanins  <= track_8_2_chanY_n15 & track_8_2_chanY_n14 & track_8_2_chanY_n11 & track_8_2_chanY_n10 & track_8_2_chanY_n7 & track_8_2_chanY_n6 & track_8_2_chanY_n3 & track_8_2_chanY_n2;
	IO_9_3_IN_pin_0_driver_mux_fanins  <= track_8_3_chanY_n13 & track_8_3_chanY_n12 & track_8_3_chanY_n9 & track_8_3_chanY_n8 & track_8_3_chanY_n5 & track_8_3_chanY_n4 & track_8_3_chanY_n1 & track_8_3_chanY_n0;
	IO_9_3_IN_pin_1_driver_mux_fanins  <= track_8_3_chanY_n15 & track_8_3_chanY_n14 & track_8_3_chanY_n11 & track_8_3_chanY_n10 & track_8_3_chanY_n7 & track_8_3_chanY_n6 & track_8_3_chanY_n3 & track_8_3_chanY_n2;
	IO_9_4_IN_pin_0_driver_mux_fanins  <= track_8_4_chanY_n13 & track_8_4_chanY_n12 & track_8_4_chanY_n9 & track_8_4_chanY_n8 & track_8_4_chanY_n5 & track_8_4_chanY_n4 & track_8_4_chanY_n1 & track_8_4_chanY_n0;
	IO_9_4_IN_pin_1_driver_mux_fanins  <= track_8_4_chanY_n15 & track_8_4_chanY_n14 & track_8_4_chanY_n11 & track_8_4_chanY_n10 & track_8_4_chanY_n7 & track_8_4_chanY_n6 & track_8_4_chanY_n3 & track_8_4_chanY_n2;
	IO_9_5_IN_pin_0_driver_mux_fanins  <= track_8_5_chanY_n13 & track_8_5_chanY_n12 & track_8_5_chanY_n9 & track_8_5_chanY_n8 & track_8_5_chanY_n5 & track_8_5_chanY_n4 & track_8_5_chanY_n1 & track_8_5_chanY_n0;
	IO_9_5_IN_pin_1_driver_mux_fanins  <= track_8_5_chanY_n15 & track_8_5_chanY_n14 & track_8_5_chanY_n11 & track_8_5_chanY_n10 & track_8_5_chanY_n7 & track_8_5_chanY_n6 & track_8_5_chanY_n3 & track_8_5_chanY_n2;
	IO_9_6_IN_pin_0_driver_mux_fanins  <= track_8_6_chanY_n13 & track_8_6_chanY_n12 & track_8_6_chanY_n9 & track_8_6_chanY_n8 & track_8_6_chanY_n5 & track_8_6_chanY_n4 & track_8_6_chanY_n1 & track_8_6_chanY_n0;
	IO_9_6_IN_pin_1_driver_mux_fanins  <= track_8_6_chanY_n15 & track_8_6_chanY_n14 & track_8_6_chanY_n11 & track_8_6_chanY_n10 & track_8_6_chanY_n7 & track_8_6_chanY_n6 & track_8_6_chanY_n3 & track_8_6_chanY_n2;

	-- Input pins selectors (selector of the mux driving the pin, i.e. the bitstream portion configuring the input pin) --
	CLB_1_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6337 downto 6336)));
	CLB_1_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6339 downto 6338)));
	CLB_1_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6341 downto 6340)));
	CLB_1_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6343 downto 6342)));
	CLB_1_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6345 downto 6344)));
	CLB_1_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6347 downto 6346)));
	CLB_1_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6349 downto 6348)));
	CLB_1_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6351 downto 6350)));
	CLB_1_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6353 downto 6352)));
	CLB_1_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6355 downto 6354)));
	CLB_1_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6357 downto 6356)));
	CLB_1_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6359 downto 6358)));
	CLB_1_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6361 downto 6360)));
	CLB_1_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6363 downto 6362)));
	CLB_1_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6365 downto 6364)));
	CLB_1_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6367 downto 6366)));
	CLB_1_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6369 downto 6368)));
	CLB_1_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6371 downto 6370)));
	CLB_1_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6373 downto 6372)));
	CLB_1_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6375 downto 6374)));
	CLB_1_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6377 downto 6376)));
	CLB_1_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6379 downto 6378)));
	CLB_1_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6381 downto 6380)));
	CLB_1_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6383 downto 6382)));
	CLB_1_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6385 downto 6384)));
	CLB_1_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6387 downto 6386)));
	CLB_1_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6389 downto 6388)));
	CLB_1_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6391 downto 6390)));
	CLB_1_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6393 downto 6392)));
	CLB_1_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6395 downto 6394)));
	CLB_1_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6397 downto 6396)));
	CLB_1_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6399 downto 6398)));
	CLB_1_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6401 downto 6400)));
	CLB_1_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6403 downto 6402)));
	CLB_1_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6405 downto 6404)));
	CLB_1_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6407 downto 6406)));
	CLB_1_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6409 downto 6408)));
	CLB_1_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6411 downto 6410)));
	CLB_1_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6413 downto 6412)));
	CLB_1_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6415 downto 6414)));
	CLB_1_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6417 downto 6416)));
	CLB_1_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6419 downto 6418)));
	CLB_1_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6421 downto 6420)));
	CLB_1_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6423 downto 6422)));
	CLB_1_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6425 downto 6424)));
	CLB_1_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6427 downto 6426)));
	CLB_1_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6429 downto 6428)));
	CLB_1_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6431 downto 6430)));
	CLB_1_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6433 downto 6432)));
	CLB_1_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6435 downto 6434)));
	CLB_1_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6437 downto 6436)));
	CLB_1_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6439 downto 6438)));
	CLB_1_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6441 downto 6440)));
	CLB_1_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6443 downto 6442)));
	CLB_1_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6445 downto 6444)));
	CLB_1_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6447 downto 6446)));
	CLB_1_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6449 downto 6448)));
	CLB_1_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6451 downto 6450)));
	CLB_1_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6453 downto 6452)));
	CLB_1_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6455 downto 6454)));
	CLB_2_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6457 downto 6456)));
	CLB_2_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6459 downto 6458)));
	CLB_2_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6461 downto 6460)));
	CLB_2_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6463 downto 6462)));
	CLB_2_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6465 downto 6464)));
	CLB_2_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6467 downto 6466)));
	CLB_2_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6469 downto 6468)));
	CLB_2_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6471 downto 6470)));
	CLB_2_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6473 downto 6472)));
	CLB_2_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6475 downto 6474)));
	CLB_2_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6477 downto 6476)));
	CLB_2_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6479 downto 6478)));
	CLB_2_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6481 downto 6480)));
	CLB_2_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6483 downto 6482)));
	CLB_2_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6485 downto 6484)));
	CLB_2_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6487 downto 6486)));
	CLB_2_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6489 downto 6488)));
	CLB_2_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6491 downto 6490)));
	CLB_2_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6493 downto 6492)));
	CLB_2_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6495 downto 6494)));
	CLB_2_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6497 downto 6496)));
	CLB_2_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6499 downto 6498)));
	CLB_2_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6501 downto 6500)));
	CLB_2_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6503 downto 6502)));
	CLB_2_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6505 downto 6504)));
	CLB_2_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6507 downto 6506)));
	CLB_2_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6509 downto 6508)));
	CLB_2_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6511 downto 6510)));
	CLB_2_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6513 downto 6512)));
	CLB_2_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6515 downto 6514)));
	CLB_2_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6517 downto 6516)));
	CLB_2_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6519 downto 6518)));
	CLB_2_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6521 downto 6520)));
	CLB_2_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6523 downto 6522)));
	CLB_2_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6525 downto 6524)));
	CLB_2_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6527 downto 6526)));
	CLB_2_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6529 downto 6528)));
	CLB_2_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6531 downto 6530)));
	CLB_2_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6533 downto 6532)));
	CLB_2_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6535 downto 6534)));
	CLB_2_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6537 downto 6536)));
	CLB_2_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6539 downto 6538)));
	CLB_2_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6541 downto 6540)));
	CLB_2_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6543 downto 6542)));
	CLB_2_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6545 downto 6544)));
	CLB_2_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6547 downto 6546)));
	CLB_2_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6549 downto 6548)));
	CLB_2_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6551 downto 6550)));
	CLB_2_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6553 downto 6552)));
	CLB_2_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6555 downto 6554)));
	CLB_2_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6557 downto 6556)));
	CLB_2_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6559 downto 6558)));
	CLB_2_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6561 downto 6560)));
	CLB_2_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6563 downto 6562)));
	CLB_2_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6565 downto 6564)));
	CLB_2_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6567 downto 6566)));
	CLB_2_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6569 downto 6568)));
	CLB_2_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6571 downto 6570)));
	CLB_2_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6573 downto 6572)));
	CLB_2_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6575 downto 6574)));
	CLB_3_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6577 downto 6576)));
	CLB_3_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6579 downto 6578)));
	CLB_3_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6581 downto 6580)));
	CLB_3_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6583 downto 6582)));
	CLB_3_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6585 downto 6584)));
	CLB_3_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6587 downto 6586)));
	CLB_3_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6589 downto 6588)));
	CLB_3_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6591 downto 6590)));
	CLB_3_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6593 downto 6592)));
	CLB_3_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6595 downto 6594)));
	CLB_3_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6597 downto 6596)));
	CLB_3_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6599 downto 6598)));
	CLB_3_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6601 downto 6600)));
	CLB_3_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6603 downto 6602)));
	CLB_3_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6605 downto 6604)));
	CLB_3_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6607 downto 6606)));
	CLB_3_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6609 downto 6608)));
	CLB_3_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6611 downto 6610)));
	CLB_3_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6613 downto 6612)));
	CLB_3_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6615 downto 6614)));
	CLB_3_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6617 downto 6616)));
	CLB_3_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6619 downto 6618)));
	CLB_3_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6621 downto 6620)));
	CLB_3_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6623 downto 6622)));
	CLB_3_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6625 downto 6624)));
	CLB_3_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6627 downto 6626)));
	CLB_3_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6629 downto 6628)));
	CLB_3_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6631 downto 6630)));
	CLB_3_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6633 downto 6632)));
	CLB_3_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6635 downto 6634)));
	CLB_3_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6637 downto 6636)));
	CLB_3_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6639 downto 6638)));
	CLB_3_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6641 downto 6640)));
	CLB_3_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6643 downto 6642)));
	CLB_3_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6645 downto 6644)));
	CLB_3_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6647 downto 6646)));
	CLB_3_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6649 downto 6648)));
	CLB_3_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6651 downto 6650)));
	CLB_3_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6653 downto 6652)));
	CLB_3_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6655 downto 6654)));
	CLB_3_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6657 downto 6656)));
	CLB_3_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6659 downto 6658)));
	CLB_3_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6661 downto 6660)));
	CLB_3_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6663 downto 6662)));
	CLB_3_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6665 downto 6664)));
	CLB_3_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6667 downto 6666)));
	CLB_3_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6669 downto 6668)));
	CLB_3_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6671 downto 6670)));
	CLB_3_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6673 downto 6672)));
	CLB_3_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6675 downto 6674)));
	CLB_3_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6677 downto 6676)));
	CLB_3_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6679 downto 6678)));
	CLB_3_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6681 downto 6680)));
	CLB_3_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6683 downto 6682)));
	CLB_3_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6685 downto 6684)));
	CLB_3_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6687 downto 6686)));
	CLB_3_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6689 downto 6688)));
	CLB_3_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6691 downto 6690)));
	CLB_3_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6693 downto 6692)));
	CLB_3_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6695 downto 6694)));
	CLB_4_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6697 downto 6696)));
	CLB_4_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6699 downto 6698)));
	CLB_4_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6701 downto 6700)));
	CLB_4_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6703 downto 6702)));
	CLB_4_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6705 downto 6704)));
	CLB_4_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6707 downto 6706)));
	CLB_4_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6709 downto 6708)));
	CLB_4_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6711 downto 6710)));
	CLB_4_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6713 downto 6712)));
	CLB_4_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6715 downto 6714)));
	CLB_4_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6717 downto 6716)));
	CLB_4_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6719 downto 6718)));
	CLB_4_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6721 downto 6720)));
	CLB_4_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6723 downto 6722)));
	CLB_4_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6725 downto 6724)));
	CLB_4_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6727 downto 6726)));
	CLB_4_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6729 downto 6728)));
	CLB_4_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6731 downto 6730)));
	CLB_4_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6733 downto 6732)));
	CLB_4_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6735 downto 6734)));
	CLB_4_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6737 downto 6736)));
	CLB_4_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6739 downto 6738)));
	CLB_4_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6741 downto 6740)));
	CLB_4_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6743 downto 6742)));
	CLB_4_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6745 downto 6744)));
	CLB_4_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6747 downto 6746)));
	CLB_4_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6749 downto 6748)));
	CLB_4_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6751 downto 6750)));
	CLB_4_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6753 downto 6752)));
	CLB_4_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6755 downto 6754)));
	CLB_4_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6757 downto 6756)));
	CLB_4_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6759 downto 6758)));
	CLB_4_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6761 downto 6760)));
	CLB_4_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6763 downto 6762)));
	CLB_4_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6765 downto 6764)));
	CLB_4_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6767 downto 6766)));
	CLB_4_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6769 downto 6768)));
	CLB_4_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6771 downto 6770)));
	CLB_4_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6773 downto 6772)));
	CLB_4_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6775 downto 6774)));
	CLB_4_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6777 downto 6776)));
	CLB_4_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6779 downto 6778)));
	CLB_4_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6781 downto 6780)));
	CLB_4_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6783 downto 6782)));
	CLB_4_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6785 downto 6784)));
	CLB_4_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6787 downto 6786)));
	CLB_4_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6789 downto 6788)));
	CLB_4_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6791 downto 6790)));
	CLB_4_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6793 downto 6792)));
	CLB_4_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6795 downto 6794)));
	CLB_4_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6797 downto 6796)));
	CLB_4_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6799 downto 6798)));
	CLB_4_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6801 downto 6800)));
	CLB_4_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6803 downto 6802)));
	CLB_4_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6805 downto 6804)));
	CLB_4_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6807 downto 6806)));
	CLB_4_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6809 downto 6808)));
	CLB_4_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6811 downto 6810)));
	CLB_4_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6813 downto 6812)));
	CLB_4_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6815 downto 6814)));
	CLB_5_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6817 downto 6816)));
	CLB_5_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6819 downto 6818)));
	CLB_5_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6821 downto 6820)));
	CLB_5_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6823 downto 6822)));
	CLB_5_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6825 downto 6824)));
	CLB_5_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6827 downto 6826)));
	CLB_5_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6829 downto 6828)));
	CLB_5_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6831 downto 6830)));
	CLB_5_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6833 downto 6832)));
	CLB_5_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6835 downto 6834)));
	CLB_5_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6837 downto 6836)));
	CLB_5_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6839 downto 6838)));
	CLB_5_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6841 downto 6840)));
	CLB_5_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6843 downto 6842)));
	CLB_5_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6845 downto 6844)));
	CLB_5_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6847 downto 6846)));
	CLB_5_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6849 downto 6848)));
	CLB_5_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6851 downto 6850)));
	CLB_5_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6853 downto 6852)));
	CLB_5_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6855 downto 6854)));
	CLB_5_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6857 downto 6856)));
	CLB_5_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6859 downto 6858)));
	CLB_5_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6861 downto 6860)));
	CLB_5_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6863 downto 6862)));
	CLB_5_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6865 downto 6864)));
	CLB_5_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6867 downto 6866)));
	CLB_5_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6869 downto 6868)));
	CLB_5_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6871 downto 6870)));
	CLB_5_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6873 downto 6872)));
	CLB_5_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6875 downto 6874)));
	CLB_5_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6877 downto 6876)));
	CLB_5_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6879 downto 6878)));
	CLB_5_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6881 downto 6880)));
	CLB_5_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6883 downto 6882)));
	CLB_5_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6885 downto 6884)));
	CLB_5_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6887 downto 6886)));
	CLB_5_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6889 downto 6888)));
	CLB_5_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6891 downto 6890)));
	CLB_5_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6893 downto 6892)));
	CLB_5_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6895 downto 6894)));
	CLB_5_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6897 downto 6896)));
	CLB_5_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6899 downto 6898)));
	CLB_5_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6901 downto 6900)));
	CLB_5_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6903 downto 6902)));
	CLB_5_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6905 downto 6904)));
	CLB_5_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6907 downto 6906)));
	CLB_5_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6909 downto 6908)));
	CLB_5_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6911 downto 6910)));
	CLB_5_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6913 downto 6912)));
	CLB_5_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6915 downto 6914)));
	CLB_5_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6917 downto 6916)));
	CLB_5_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6919 downto 6918)));
	CLB_5_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6921 downto 6920)));
	CLB_5_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6923 downto 6922)));
	CLB_5_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6925 downto 6924)));
	CLB_5_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6927 downto 6926)));
	CLB_5_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6929 downto 6928)));
	CLB_5_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6931 downto 6930)));
	CLB_5_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6933 downto 6932)));
	CLB_5_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6935 downto 6934)));
	CLB_6_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6937 downto 6936)));
	CLB_6_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6939 downto 6938)));
	CLB_6_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6941 downto 6940)));
	CLB_6_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6943 downto 6942)));
	CLB_6_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6945 downto 6944)));
	CLB_6_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6947 downto 6946)));
	CLB_6_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6949 downto 6948)));
	CLB_6_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6951 downto 6950)));
	CLB_6_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6953 downto 6952)));
	CLB_6_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6955 downto 6954)));
	CLB_6_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6957 downto 6956)));
	CLB_6_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6959 downto 6958)));
	CLB_6_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6961 downto 6960)));
	CLB_6_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6963 downto 6962)));
	CLB_6_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6965 downto 6964)));
	CLB_6_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6967 downto 6966)));
	CLB_6_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6969 downto 6968)));
	CLB_6_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6971 downto 6970)));
	CLB_6_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6973 downto 6972)));
	CLB_6_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6975 downto 6974)));
	CLB_6_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6977 downto 6976)));
	CLB_6_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6979 downto 6978)));
	CLB_6_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(6981 downto 6980)));
	CLB_6_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(6983 downto 6982)));
	CLB_6_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(6985 downto 6984)));
	CLB_6_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(6987 downto 6986)));
	CLB_6_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(6989 downto 6988)));
	CLB_6_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(6991 downto 6990)));
	CLB_6_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(6993 downto 6992)));
	CLB_6_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(6995 downto 6994)));
	CLB_6_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(6997 downto 6996)));
	CLB_6_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(6999 downto 6998)));
	CLB_6_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7001 downto 7000)));
	CLB_6_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7003 downto 7002)));
	CLB_6_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7005 downto 7004)));
	CLB_6_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7007 downto 7006)));
	CLB_6_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7009 downto 7008)));
	CLB_6_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7011 downto 7010)));
	CLB_6_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7013 downto 7012)));
	CLB_6_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7015 downto 7014)));
	CLB_6_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7017 downto 7016)));
	CLB_6_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7019 downto 7018)));
	CLB_6_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7021 downto 7020)));
	CLB_6_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7023 downto 7022)));
	CLB_6_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7025 downto 7024)));
	CLB_6_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7027 downto 7026)));
	CLB_6_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7029 downto 7028)));
	CLB_6_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7031 downto 7030)));
	CLB_6_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7033 downto 7032)));
	CLB_6_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7035 downto 7034)));
	CLB_6_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7037 downto 7036)));
	CLB_6_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7039 downto 7038)));
	CLB_6_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7041 downto 7040)));
	CLB_6_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7043 downto 7042)));
	CLB_6_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7045 downto 7044)));
	CLB_6_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7047 downto 7046)));
	CLB_6_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7049 downto 7048)));
	CLB_6_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7051 downto 7050)));
	CLB_6_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7053 downto 7052)));
	CLB_6_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7055 downto 7054)));
	CLB_7_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7057 downto 7056)));
	CLB_7_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7059 downto 7058)));
	CLB_7_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7061 downto 7060)));
	CLB_7_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7063 downto 7062)));
	CLB_7_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7065 downto 7064)));
	CLB_7_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7067 downto 7066)));
	CLB_7_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7069 downto 7068)));
	CLB_7_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7071 downto 7070)));
	CLB_7_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7073 downto 7072)));
	CLB_7_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7075 downto 7074)));
	CLB_7_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7077 downto 7076)));
	CLB_7_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7079 downto 7078)));
	CLB_7_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7081 downto 7080)));
	CLB_7_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7083 downto 7082)));
	CLB_7_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7085 downto 7084)));
	CLB_7_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7087 downto 7086)));
	CLB_7_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7089 downto 7088)));
	CLB_7_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7091 downto 7090)));
	CLB_7_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7093 downto 7092)));
	CLB_7_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7095 downto 7094)));
	CLB_7_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7097 downto 7096)));
	CLB_7_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7099 downto 7098)));
	CLB_7_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7101 downto 7100)));
	CLB_7_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7103 downto 7102)));
	CLB_7_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7105 downto 7104)));
	CLB_7_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7107 downto 7106)));
	CLB_7_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7109 downto 7108)));
	CLB_7_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7111 downto 7110)));
	CLB_7_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7113 downto 7112)));
	CLB_7_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7115 downto 7114)));
	CLB_7_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7117 downto 7116)));
	CLB_7_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7119 downto 7118)));
	CLB_7_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7121 downto 7120)));
	CLB_7_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7123 downto 7122)));
	CLB_7_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7125 downto 7124)));
	CLB_7_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7127 downto 7126)));
	CLB_7_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7129 downto 7128)));
	CLB_7_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7131 downto 7130)));
	CLB_7_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7133 downto 7132)));
	CLB_7_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7135 downto 7134)));
	CLB_7_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7137 downto 7136)));
	CLB_7_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7139 downto 7138)));
	CLB_7_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7141 downto 7140)));
	CLB_7_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7143 downto 7142)));
	CLB_7_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7145 downto 7144)));
	CLB_7_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7147 downto 7146)));
	CLB_7_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7149 downto 7148)));
	CLB_7_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7151 downto 7150)));
	CLB_7_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7153 downto 7152)));
	CLB_7_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7155 downto 7154)));
	CLB_7_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7157 downto 7156)));
	CLB_7_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7159 downto 7158)));
	CLB_7_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7161 downto 7160)));
	CLB_7_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7163 downto 7162)));
	CLB_7_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7165 downto 7164)));
	CLB_7_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7167 downto 7166)));
	CLB_7_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7169 downto 7168)));
	CLB_7_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7171 downto 7170)));
	CLB_7_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7173 downto 7172)));
	CLB_7_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7175 downto 7174)));
	CLB_8_1_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7177 downto 7176)));
	CLB_8_1_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7179 downto 7178)));
	CLB_8_1_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7181 downto 7180)));
	CLB_8_1_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7183 downto 7182)));
	CLB_8_1_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7185 downto 7184)));
	CLB_8_1_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7187 downto 7186)));
	CLB_8_1_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7189 downto 7188)));
	CLB_8_1_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7191 downto 7190)));
	CLB_8_1_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7193 downto 7192)));
	CLB_8_1_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7195 downto 7194)));
	CLB_8_2_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7197 downto 7196)));
	CLB_8_2_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7199 downto 7198)));
	CLB_8_2_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7201 downto 7200)));
	CLB_8_2_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7203 downto 7202)));
	CLB_8_2_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7205 downto 7204)));
	CLB_8_2_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7207 downto 7206)));
	CLB_8_2_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7209 downto 7208)));
	CLB_8_2_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7211 downto 7210)));
	CLB_8_2_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7213 downto 7212)));
	CLB_8_2_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7215 downto 7214)));
	CLB_8_3_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7217 downto 7216)));
	CLB_8_3_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7219 downto 7218)));
	CLB_8_3_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7221 downto 7220)));
	CLB_8_3_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7223 downto 7222)));
	CLB_8_3_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7225 downto 7224)));
	CLB_8_3_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7227 downto 7226)));
	CLB_8_3_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7229 downto 7228)));
	CLB_8_3_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7231 downto 7230)));
	CLB_8_3_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7233 downto 7232)));
	CLB_8_3_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7235 downto 7234)));
	CLB_8_4_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7237 downto 7236)));
	CLB_8_4_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7239 downto 7238)));
	CLB_8_4_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7241 downto 7240)));
	CLB_8_4_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7243 downto 7242)));
	CLB_8_4_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7245 downto 7244)));
	CLB_8_4_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7247 downto 7246)));
	CLB_8_4_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7249 downto 7248)));
	CLB_8_4_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7251 downto 7250)));
	CLB_8_4_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7253 downto 7252)));
	CLB_8_4_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7255 downto 7254)));
	CLB_8_5_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7257 downto 7256)));
	CLB_8_5_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7259 downto 7258)));
	CLB_8_5_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7261 downto 7260)));
	CLB_8_5_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7263 downto 7262)));
	CLB_8_5_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7265 downto 7264)));
	CLB_8_5_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7267 downto 7266)));
	CLB_8_5_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7269 downto 7268)));
	CLB_8_5_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7271 downto 7270)));
	CLB_8_5_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7273 downto 7272)));
	CLB_8_5_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7275 downto 7274)));
	CLB_8_6_IN_pin_0_driver_mux_selector <= to_integer(unsigned(config(7277 downto 7276)));
	CLB_8_6_IN_pin_1_driver_mux_selector <= to_integer(unsigned(config(7279 downto 7278)));
	CLB_8_6_IN_pin_2_driver_mux_selector <= to_integer(unsigned(config(7281 downto 7280)));
	CLB_8_6_IN_pin_3_driver_mux_selector <= to_integer(unsigned(config(7283 downto 7282)));
	CLB_8_6_IN_pin_4_driver_mux_selector <= to_integer(unsigned(config(7285 downto 7284)));
	CLB_8_6_IN_pin_5_driver_mux_selector <= to_integer(unsigned(config(7287 downto 7286)));
	CLB_8_6_IN_pin_6_driver_mux_selector <= to_integer(unsigned(config(7289 downto 7288)));
	CLB_8_6_IN_pin_7_driver_mux_selector <= to_integer(unsigned(config(7291 downto 7290)));
	CLB_8_6_IN_pin_8_driver_mux_selector <= to_integer(unsigned(config(7293 downto 7292)));
	CLB_8_6_IN_pin_9_driver_mux_selector <= to_integer(unsigned(config(7295 downto 7294)));
	IO_0_1_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7298 downto 7296)));
	IO_0_1_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7301 downto 7299)));
	IO_0_2_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7304 downto 7302)));
	IO_0_2_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7307 downto 7305)));
	IO_0_3_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7310 downto 7308)));
	IO_0_3_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7313 downto 7311)));
	IO_0_4_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7316 downto 7314)));
	IO_0_4_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7319 downto 7317)));
	IO_0_5_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7322 downto 7320)));
	IO_0_5_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7325 downto 7323)));
	IO_0_6_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7328 downto 7326)));
	IO_0_6_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7331 downto 7329)));
	IO_1_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7334 downto 7332)));
	IO_1_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7337 downto 7335)));
	IO_1_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7340 downto 7338)));
	IO_1_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7343 downto 7341)));
	IO_2_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7346 downto 7344)));
	IO_2_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7349 downto 7347)));
	IO_2_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7352 downto 7350)));
	IO_2_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7355 downto 7353)));
	IO_3_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7358 downto 7356)));
	IO_3_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7361 downto 7359)));
	IO_3_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7364 downto 7362)));
	IO_3_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7367 downto 7365)));
	IO_4_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7370 downto 7368)));
	IO_4_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7373 downto 7371)));
	IO_4_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7376 downto 7374)));
	IO_4_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7379 downto 7377)));
	IO_5_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7382 downto 7380)));
	IO_5_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7385 downto 7383)));
	IO_5_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7388 downto 7386)));
	IO_5_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7391 downto 7389)));
	IO_6_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7394 downto 7392)));
	IO_6_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7397 downto 7395)));
	IO_6_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7400 downto 7398)));
	IO_6_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7403 downto 7401)));
	IO_7_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7406 downto 7404)));
	IO_7_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7409 downto 7407)));
	IO_7_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7412 downto 7410)));
	IO_7_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7415 downto 7413)));
	IO_8_0_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7418 downto 7416)));
	IO_8_0_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7421 downto 7419)));
	IO_8_7_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7424 downto 7422)));
	IO_8_7_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7427 downto 7425)));
	IO_9_1_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7430 downto 7428)));
	IO_9_1_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7433 downto 7431)));
	IO_9_2_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7436 downto 7434)));
	IO_9_2_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7439 downto 7437)));
	IO_9_3_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7442 downto 7440)));
	IO_9_3_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7445 downto 7443)));
	IO_9_4_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7448 downto 7446)));
	IO_9_4_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7451 downto 7449)));
	IO_9_5_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7454 downto 7452)));
	IO_9_5_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7457 downto 7455)));
	IO_9_6_IN_pin_0_driver_mux_selector  <= to_integer(unsigned(config(7460 downto 7458)));
	IO_9_6_IN_pin_1_driver_mux_selector  <= to_integer(unsigned(config(7463 downto 7461)));

	-- Input pins (for CLBs and IOs) --
	CLB_1_1_IN_pin_0 <= CLB_1_1_IN_pin_0_driver_mux_fanins(CLB_1_1_IN_pin_0_driver_mux_selector);
	CLB_1_1_IN_pin_1 <= CLB_1_1_IN_pin_1_driver_mux_fanins(CLB_1_1_IN_pin_1_driver_mux_selector);
	CLB_1_1_IN_pin_2 <= CLB_1_1_IN_pin_2_driver_mux_fanins(CLB_1_1_IN_pin_2_driver_mux_selector);
	CLB_1_1_IN_pin_3 <= CLB_1_1_IN_pin_3_driver_mux_fanins(CLB_1_1_IN_pin_3_driver_mux_selector);
	CLB_1_1_IN_pin_4 <= CLB_1_1_IN_pin_4_driver_mux_fanins(CLB_1_1_IN_pin_4_driver_mux_selector);
	CLB_1_1_IN_pin_5 <= CLB_1_1_IN_pin_5_driver_mux_fanins(CLB_1_1_IN_pin_5_driver_mux_selector);
	CLB_1_1_IN_pin_6 <= CLB_1_1_IN_pin_6_driver_mux_fanins(CLB_1_1_IN_pin_6_driver_mux_selector);
	CLB_1_1_IN_pin_7 <= CLB_1_1_IN_pin_7_driver_mux_fanins(CLB_1_1_IN_pin_7_driver_mux_selector);
	CLB_1_1_IN_pin_8 <= CLB_1_1_IN_pin_8_driver_mux_fanins(CLB_1_1_IN_pin_8_driver_mux_selector);
	CLB_1_1_IN_pin_9 <= CLB_1_1_IN_pin_9_driver_mux_fanins(CLB_1_1_IN_pin_9_driver_mux_selector);
	CLB_1_2_IN_pin_0 <= CLB_1_2_IN_pin_0_driver_mux_fanins(CLB_1_2_IN_pin_0_driver_mux_selector);
	CLB_1_2_IN_pin_1 <= CLB_1_2_IN_pin_1_driver_mux_fanins(CLB_1_2_IN_pin_1_driver_mux_selector);
	CLB_1_2_IN_pin_2 <= CLB_1_2_IN_pin_2_driver_mux_fanins(CLB_1_2_IN_pin_2_driver_mux_selector);
	CLB_1_2_IN_pin_3 <= CLB_1_2_IN_pin_3_driver_mux_fanins(CLB_1_2_IN_pin_3_driver_mux_selector);
	CLB_1_2_IN_pin_4 <= CLB_1_2_IN_pin_4_driver_mux_fanins(CLB_1_2_IN_pin_4_driver_mux_selector);
	CLB_1_2_IN_pin_5 <= CLB_1_2_IN_pin_5_driver_mux_fanins(CLB_1_2_IN_pin_5_driver_mux_selector);
	CLB_1_2_IN_pin_6 <= CLB_1_2_IN_pin_6_driver_mux_fanins(CLB_1_2_IN_pin_6_driver_mux_selector);
	CLB_1_2_IN_pin_7 <= CLB_1_2_IN_pin_7_driver_mux_fanins(CLB_1_2_IN_pin_7_driver_mux_selector);
	CLB_1_2_IN_pin_8 <= CLB_1_2_IN_pin_8_driver_mux_fanins(CLB_1_2_IN_pin_8_driver_mux_selector);
	CLB_1_2_IN_pin_9 <= CLB_1_2_IN_pin_9_driver_mux_fanins(CLB_1_2_IN_pin_9_driver_mux_selector);
	CLB_1_3_IN_pin_0 <= CLB_1_3_IN_pin_0_driver_mux_fanins(CLB_1_3_IN_pin_0_driver_mux_selector);
	CLB_1_3_IN_pin_1 <= CLB_1_3_IN_pin_1_driver_mux_fanins(CLB_1_3_IN_pin_1_driver_mux_selector);
	CLB_1_3_IN_pin_2 <= CLB_1_3_IN_pin_2_driver_mux_fanins(CLB_1_3_IN_pin_2_driver_mux_selector);
	CLB_1_3_IN_pin_3 <= CLB_1_3_IN_pin_3_driver_mux_fanins(CLB_1_3_IN_pin_3_driver_mux_selector);
	CLB_1_3_IN_pin_4 <= CLB_1_3_IN_pin_4_driver_mux_fanins(CLB_1_3_IN_pin_4_driver_mux_selector);
	CLB_1_3_IN_pin_5 <= CLB_1_3_IN_pin_5_driver_mux_fanins(CLB_1_3_IN_pin_5_driver_mux_selector);
	CLB_1_3_IN_pin_6 <= CLB_1_3_IN_pin_6_driver_mux_fanins(CLB_1_3_IN_pin_6_driver_mux_selector);
	CLB_1_3_IN_pin_7 <= CLB_1_3_IN_pin_7_driver_mux_fanins(CLB_1_3_IN_pin_7_driver_mux_selector);
	CLB_1_3_IN_pin_8 <= CLB_1_3_IN_pin_8_driver_mux_fanins(CLB_1_3_IN_pin_8_driver_mux_selector);
	CLB_1_3_IN_pin_9 <= CLB_1_3_IN_pin_9_driver_mux_fanins(CLB_1_3_IN_pin_9_driver_mux_selector);
	CLB_1_4_IN_pin_0 <= CLB_1_4_IN_pin_0_driver_mux_fanins(CLB_1_4_IN_pin_0_driver_mux_selector);
	CLB_1_4_IN_pin_1 <= CLB_1_4_IN_pin_1_driver_mux_fanins(CLB_1_4_IN_pin_1_driver_mux_selector);
	CLB_1_4_IN_pin_2 <= CLB_1_4_IN_pin_2_driver_mux_fanins(CLB_1_4_IN_pin_2_driver_mux_selector);
	CLB_1_4_IN_pin_3 <= CLB_1_4_IN_pin_3_driver_mux_fanins(CLB_1_4_IN_pin_3_driver_mux_selector);
	CLB_1_4_IN_pin_4 <= CLB_1_4_IN_pin_4_driver_mux_fanins(CLB_1_4_IN_pin_4_driver_mux_selector);
	CLB_1_4_IN_pin_5 <= CLB_1_4_IN_pin_5_driver_mux_fanins(CLB_1_4_IN_pin_5_driver_mux_selector);
	CLB_1_4_IN_pin_6 <= CLB_1_4_IN_pin_6_driver_mux_fanins(CLB_1_4_IN_pin_6_driver_mux_selector);
	CLB_1_4_IN_pin_7 <= CLB_1_4_IN_pin_7_driver_mux_fanins(CLB_1_4_IN_pin_7_driver_mux_selector);
	CLB_1_4_IN_pin_8 <= CLB_1_4_IN_pin_8_driver_mux_fanins(CLB_1_4_IN_pin_8_driver_mux_selector);
	CLB_1_4_IN_pin_9 <= CLB_1_4_IN_pin_9_driver_mux_fanins(CLB_1_4_IN_pin_9_driver_mux_selector);
	CLB_1_5_IN_pin_0 <= CLB_1_5_IN_pin_0_driver_mux_fanins(CLB_1_5_IN_pin_0_driver_mux_selector);
	CLB_1_5_IN_pin_1 <= CLB_1_5_IN_pin_1_driver_mux_fanins(CLB_1_5_IN_pin_1_driver_mux_selector);
	CLB_1_5_IN_pin_2 <= CLB_1_5_IN_pin_2_driver_mux_fanins(CLB_1_5_IN_pin_2_driver_mux_selector);
	CLB_1_5_IN_pin_3 <= CLB_1_5_IN_pin_3_driver_mux_fanins(CLB_1_5_IN_pin_3_driver_mux_selector);
	CLB_1_5_IN_pin_4 <= CLB_1_5_IN_pin_4_driver_mux_fanins(CLB_1_5_IN_pin_4_driver_mux_selector);
	CLB_1_5_IN_pin_5 <= CLB_1_5_IN_pin_5_driver_mux_fanins(CLB_1_5_IN_pin_5_driver_mux_selector);
	CLB_1_5_IN_pin_6 <= CLB_1_5_IN_pin_6_driver_mux_fanins(CLB_1_5_IN_pin_6_driver_mux_selector);
	CLB_1_5_IN_pin_7 <= CLB_1_5_IN_pin_7_driver_mux_fanins(CLB_1_5_IN_pin_7_driver_mux_selector);
	CLB_1_5_IN_pin_8 <= CLB_1_5_IN_pin_8_driver_mux_fanins(CLB_1_5_IN_pin_8_driver_mux_selector);
	CLB_1_5_IN_pin_9 <= CLB_1_5_IN_pin_9_driver_mux_fanins(CLB_1_5_IN_pin_9_driver_mux_selector);
	CLB_1_6_IN_pin_0 <= CLB_1_6_IN_pin_0_driver_mux_fanins(CLB_1_6_IN_pin_0_driver_mux_selector);
	CLB_1_6_IN_pin_1 <= CLB_1_6_IN_pin_1_driver_mux_fanins(CLB_1_6_IN_pin_1_driver_mux_selector);
	CLB_1_6_IN_pin_2 <= CLB_1_6_IN_pin_2_driver_mux_fanins(CLB_1_6_IN_pin_2_driver_mux_selector);
	CLB_1_6_IN_pin_3 <= CLB_1_6_IN_pin_3_driver_mux_fanins(CLB_1_6_IN_pin_3_driver_mux_selector);
	CLB_1_6_IN_pin_4 <= CLB_1_6_IN_pin_4_driver_mux_fanins(CLB_1_6_IN_pin_4_driver_mux_selector);
	CLB_1_6_IN_pin_5 <= CLB_1_6_IN_pin_5_driver_mux_fanins(CLB_1_6_IN_pin_5_driver_mux_selector);
	CLB_1_6_IN_pin_6 <= CLB_1_6_IN_pin_6_driver_mux_fanins(CLB_1_6_IN_pin_6_driver_mux_selector);
	CLB_1_6_IN_pin_7 <= CLB_1_6_IN_pin_7_driver_mux_fanins(CLB_1_6_IN_pin_7_driver_mux_selector);
	CLB_1_6_IN_pin_8 <= CLB_1_6_IN_pin_8_driver_mux_fanins(CLB_1_6_IN_pin_8_driver_mux_selector);
	CLB_1_6_IN_pin_9 <= CLB_1_6_IN_pin_9_driver_mux_fanins(CLB_1_6_IN_pin_9_driver_mux_selector);
	CLB_2_1_IN_pin_0 <= CLB_2_1_IN_pin_0_driver_mux_fanins(CLB_2_1_IN_pin_0_driver_mux_selector);
	CLB_2_1_IN_pin_1 <= CLB_2_1_IN_pin_1_driver_mux_fanins(CLB_2_1_IN_pin_1_driver_mux_selector);
	CLB_2_1_IN_pin_2 <= CLB_2_1_IN_pin_2_driver_mux_fanins(CLB_2_1_IN_pin_2_driver_mux_selector);
	CLB_2_1_IN_pin_3 <= CLB_2_1_IN_pin_3_driver_mux_fanins(CLB_2_1_IN_pin_3_driver_mux_selector);
	CLB_2_1_IN_pin_4 <= CLB_2_1_IN_pin_4_driver_mux_fanins(CLB_2_1_IN_pin_4_driver_mux_selector);
	CLB_2_1_IN_pin_5 <= CLB_2_1_IN_pin_5_driver_mux_fanins(CLB_2_1_IN_pin_5_driver_mux_selector);
	CLB_2_1_IN_pin_6 <= CLB_2_1_IN_pin_6_driver_mux_fanins(CLB_2_1_IN_pin_6_driver_mux_selector);
	CLB_2_1_IN_pin_7 <= CLB_2_1_IN_pin_7_driver_mux_fanins(CLB_2_1_IN_pin_7_driver_mux_selector);
	CLB_2_1_IN_pin_8 <= CLB_2_1_IN_pin_8_driver_mux_fanins(CLB_2_1_IN_pin_8_driver_mux_selector);
	CLB_2_1_IN_pin_9 <= CLB_2_1_IN_pin_9_driver_mux_fanins(CLB_2_1_IN_pin_9_driver_mux_selector);
	CLB_2_2_IN_pin_0 <= CLB_2_2_IN_pin_0_driver_mux_fanins(CLB_2_2_IN_pin_0_driver_mux_selector);
	CLB_2_2_IN_pin_1 <= CLB_2_2_IN_pin_1_driver_mux_fanins(CLB_2_2_IN_pin_1_driver_mux_selector);
	CLB_2_2_IN_pin_2 <= CLB_2_2_IN_pin_2_driver_mux_fanins(CLB_2_2_IN_pin_2_driver_mux_selector);
	CLB_2_2_IN_pin_3 <= CLB_2_2_IN_pin_3_driver_mux_fanins(CLB_2_2_IN_pin_3_driver_mux_selector);
	CLB_2_2_IN_pin_4 <= CLB_2_2_IN_pin_4_driver_mux_fanins(CLB_2_2_IN_pin_4_driver_mux_selector);
	CLB_2_2_IN_pin_5 <= CLB_2_2_IN_pin_5_driver_mux_fanins(CLB_2_2_IN_pin_5_driver_mux_selector);
	CLB_2_2_IN_pin_6 <= CLB_2_2_IN_pin_6_driver_mux_fanins(CLB_2_2_IN_pin_6_driver_mux_selector);
	CLB_2_2_IN_pin_7 <= CLB_2_2_IN_pin_7_driver_mux_fanins(CLB_2_2_IN_pin_7_driver_mux_selector);
	CLB_2_2_IN_pin_8 <= CLB_2_2_IN_pin_8_driver_mux_fanins(CLB_2_2_IN_pin_8_driver_mux_selector);
	CLB_2_2_IN_pin_9 <= CLB_2_2_IN_pin_9_driver_mux_fanins(CLB_2_2_IN_pin_9_driver_mux_selector);
	CLB_2_3_IN_pin_0 <= CLB_2_3_IN_pin_0_driver_mux_fanins(CLB_2_3_IN_pin_0_driver_mux_selector);
	CLB_2_3_IN_pin_1 <= CLB_2_3_IN_pin_1_driver_mux_fanins(CLB_2_3_IN_pin_1_driver_mux_selector);
	CLB_2_3_IN_pin_2 <= CLB_2_3_IN_pin_2_driver_mux_fanins(CLB_2_3_IN_pin_2_driver_mux_selector);
	CLB_2_3_IN_pin_3 <= CLB_2_3_IN_pin_3_driver_mux_fanins(CLB_2_3_IN_pin_3_driver_mux_selector);
	CLB_2_3_IN_pin_4 <= CLB_2_3_IN_pin_4_driver_mux_fanins(CLB_2_3_IN_pin_4_driver_mux_selector);
	CLB_2_3_IN_pin_5 <= CLB_2_3_IN_pin_5_driver_mux_fanins(CLB_2_3_IN_pin_5_driver_mux_selector);
	CLB_2_3_IN_pin_6 <= CLB_2_3_IN_pin_6_driver_mux_fanins(CLB_2_3_IN_pin_6_driver_mux_selector);
	CLB_2_3_IN_pin_7 <= CLB_2_3_IN_pin_7_driver_mux_fanins(CLB_2_3_IN_pin_7_driver_mux_selector);
	CLB_2_3_IN_pin_8 <= CLB_2_3_IN_pin_8_driver_mux_fanins(CLB_2_3_IN_pin_8_driver_mux_selector);
	CLB_2_3_IN_pin_9 <= CLB_2_3_IN_pin_9_driver_mux_fanins(CLB_2_3_IN_pin_9_driver_mux_selector);
	CLB_2_4_IN_pin_0 <= CLB_2_4_IN_pin_0_driver_mux_fanins(CLB_2_4_IN_pin_0_driver_mux_selector);
	CLB_2_4_IN_pin_1 <= CLB_2_4_IN_pin_1_driver_mux_fanins(CLB_2_4_IN_pin_1_driver_mux_selector);
	CLB_2_4_IN_pin_2 <= CLB_2_4_IN_pin_2_driver_mux_fanins(CLB_2_4_IN_pin_2_driver_mux_selector);
	CLB_2_4_IN_pin_3 <= CLB_2_4_IN_pin_3_driver_mux_fanins(CLB_2_4_IN_pin_3_driver_mux_selector);
	CLB_2_4_IN_pin_4 <= CLB_2_4_IN_pin_4_driver_mux_fanins(CLB_2_4_IN_pin_4_driver_mux_selector);
	CLB_2_4_IN_pin_5 <= CLB_2_4_IN_pin_5_driver_mux_fanins(CLB_2_4_IN_pin_5_driver_mux_selector);
	CLB_2_4_IN_pin_6 <= CLB_2_4_IN_pin_6_driver_mux_fanins(CLB_2_4_IN_pin_6_driver_mux_selector);
	CLB_2_4_IN_pin_7 <= CLB_2_4_IN_pin_7_driver_mux_fanins(CLB_2_4_IN_pin_7_driver_mux_selector);
	CLB_2_4_IN_pin_8 <= CLB_2_4_IN_pin_8_driver_mux_fanins(CLB_2_4_IN_pin_8_driver_mux_selector);
	CLB_2_4_IN_pin_9 <= CLB_2_4_IN_pin_9_driver_mux_fanins(CLB_2_4_IN_pin_9_driver_mux_selector);
	CLB_2_5_IN_pin_0 <= CLB_2_5_IN_pin_0_driver_mux_fanins(CLB_2_5_IN_pin_0_driver_mux_selector);
	CLB_2_5_IN_pin_1 <= CLB_2_5_IN_pin_1_driver_mux_fanins(CLB_2_5_IN_pin_1_driver_mux_selector);
	CLB_2_5_IN_pin_2 <= CLB_2_5_IN_pin_2_driver_mux_fanins(CLB_2_5_IN_pin_2_driver_mux_selector);
	CLB_2_5_IN_pin_3 <= CLB_2_5_IN_pin_3_driver_mux_fanins(CLB_2_5_IN_pin_3_driver_mux_selector);
	CLB_2_5_IN_pin_4 <= CLB_2_5_IN_pin_4_driver_mux_fanins(CLB_2_5_IN_pin_4_driver_mux_selector);
	CLB_2_5_IN_pin_5 <= CLB_2_5_IN_pin_5_driver_mux_fanins(CLB_2_5_IN_pin_5_driver_mux_selector);
	CLB_2_5_IN_pin_6 <= CLB_2_5_IN_pin_6_driver_mux_fanins(CLB_2_5_IN_pin_6_driver_mux_selector);
	CLB_2_5_IN_pin_7 <= CLB_2_5_IN_pin_7_driver_mux_fanins(CLB_2_5_IN_pin_7_driver_mux_selector);
	CLB_2_5_IN_pin_8 <= CLB_2_5_IN_pin_8_driver_mux_fanins(CLB_2_5_IN_pin_8_driver_mux_selector);
	CLB_2_5_IN_pin_9 <= CLB_2_5_IN_pin_9_driver_mux_fanins(CLB_2_5_IN_pin_9_driver_mux_selector);
	CLB_2_6_IN_pin_0 <= CLB_2_6_IN_pin_0_driver_mux_fanins(CLB_2_6_IN_pin_0_driver_mux_selector);
	CLB_2_6_IN_pin_1 <= CLB_2_6_IN_pin_1_driver_mux_fanins(CLB_2_6_IN_pin_1_driver_mux_selector);
	CLB_2_6_IN_pin_2 <= CLB_2_6_IN_pin_2_driver_mux_fanins(CLB_2_6_IN_pin_2_driver_mux_selector);
	CLB_2_6_IN_pin_3 <= CLB_2_6_IN_pin_3_driver_mux_fanins(CLB_2_6_IN_pin_3_driver_mux_selector);
	CLB_2_6_IN_pin_4 <= CLB_2_6_IN_pin_4_driver_mux_fanins(CLB_2_6_IN_pin_4_driver_mux_selector);
	CLB_2_6_IN_pin_5 <= CLB_2_6_IN_pin_5_driver_mux_fanins(CLB_2_6_IN_pin_5_driver_mux_selector);
	CLB_2_6_IN_pin_6 <= CLB_2_6_IN_pin_6_driver_mux_fanins(CLB_2_6_IN_pin_6_driver_mux_selector);
	CLB_2_6_IN_pin_7 <= CLB_2_6_IN_pin_7_driver_mux_fanins(CLB_2_6_IN_pin_7_driver_mux_selector);
	CLB_2_6_IN_pin_8 <= CLB_2_6_IN_pin_8_driver_mux_fanins(CLB_2_6_IN_pin_8_driver_mux_selector);
	CLB_2_6_IN_pin_9 <= CLB_2_6_IN_pin_9_driver_mux_fanins(CLB_2_6_IN_pin_9_driver_mux_selector);
	CLB_3_1_IN_pin_0 <= CLB_3_1_IN_pin_0_driver_mux_fanins(CLB_3_1_IN_pin_0_driver_mux_selector);
	CLB_3_1_IN_pin_1 <= CLB_3_1_IN_pin_1_driver_mux_fanins(CLB_3_1_IN_pin_1_driver_mux_selector);
	CLB_3_1_IN_pin_2 <= CLB_3_1_IN_pin_2_driver_mux_fanins(CLB_3_1_IN_pin_2_driver_mux_selector);
	CLB_3_1_IN_pin_3 <= CLB_3_1_IN_pin_3_driver_mux_fanins(CLB_3_1_IN_pin_3_driver_mux_selector);
	CLB_3_1_IN_pin_4 <= CLB_3_1_IN_pin_4_driver_mux_fanins(CLB_3_1_IN_pin_4_driver_mux_selector);
	CLB_3_1_IN_pin_5 <= CLB_3_1_IN_pin_5_driver_mux_fanins(CLB_3_1_IN_pin_5_driver_mux_selector);
	CLB_3_1_IN_pin_6 <= CLB_3_1_IN_pin_6_driver_mux_fanins(CLB_3_1_IN_pin_6_driver_mux_selector);
	CLB_3_1_IN_pin_7 <= CLB_3_1_IN_pin_7_driver_mux_fanins(CLB_3_1_IN_pin_7_driver_mux_selector);
	CLB_3_1_IN_pin_8 <= CLB_3_1_IN_pin_8_driver_mux_fanins(CLB_3_1_IN_pin_8_driver_mux_selector);
	CLB_3_1_IN_pin_9 <= CLB_3_1_IN_pin_9_driver_mux_fanins(CLB_3_1_IN_pin_9_driver_mux_selector);
	CLB_3_2_IN_pin_0 <= CLB_3_2_IN_pin_0_driver_mux_fanins(CLB_3_2_IN_pin_0_driver_mux_selector);
	CLB_3_2_IN_pin_1 <= CLB_3_2_IN_pin_1_driver_mux_fanins(CLB_3_2_IN_pin_1_driver_mux_selector);
	CLB_3_2_IN_pin_2 <= CLB_3_2_IN_pin_2_driver_mux_fanins(CLB_3_2_IN_pin_2_driver_mux_selector);
	CLB_3_2_IN_pin_3 <= CLB_3_2_IN_pin_3_driver_mux_fanins(CLB_3_2_IN_pin_3_driver_mux_selector);
	CLB_3_2_IN_pin_4 <= CLB_3_2_IN_pin_4_driver_mux_fanins(CLB_3_2_IN_pin_4_driver_mux_selector);
	CLB_3_2_IN_pin_5 <= CLB_3_2_IN_pin_5_driver_mux_fanins(CLB_3_2_IN_pin_5_driver_mux_selector);
	CLB_3_2_IN_pin_6 <= CLB_3_2_IN_pin_6_driver_mux_fanins(CLB_3_2_IN_pin_6_driver_mux_selector);
	CLB_3_2_IN_pin_7 <= CLB_3_2_IN_pin_7_driver_mux_fanins(CLB_3_2_IN_pin_7_driver_mux_selector);
	CLB_3_2_IN_pin_8 <= CLB_3_2_IN_pin_8_driver_mux_fanins(CLB_3_2_IN_pin_8_driver_mux_selector);
	CLB_3_2_IN_pin_9 <= CLB_3_2_IN_pin_9_driver_mux_fanins(CLB_3_2_IN_pin_9_driver_mux_selector);
	CLB_3_3_IN_pin_0 <= CLB_3_3_IN_pin_0_driver_mux_fanins(CLB_3_3_IN_pin_0_driver_mux_selector);
	CLB_3_3_IN_pin_1 <= CLB_3_3_IN_pin_1_driver_mux_fanins(CLB_3_3_IN_pin_1_driver_mux_selector);
	CLB_3_3_IN_pin_2 <= CLB_3_3_IN_pin_2_driver_mux_fanins(CLB_3_3_IN_pin_2_driver_mux_selector);
	CLB_3_3_IN_pin_3 <= CLB_3_3_IN_pin_3_driver_mux_fanins(CLB_3_3_IN_pin_3_driver_mux_selector);
	CLB_3_3_IN_pin_4 <= CLB_3_3_IN_pin_4_driver_mux_fanins(CLB_3_3_IN_pin_4_driver_mux_selector);
	CLB_3_3_IN_pin_5 <= CLB_3_3_IN_pin_5_driver_mux_fanins(CLB_3_3_IN_pin_5_driver_mux_selector);
	CLB_3_3_IN_pin_6 <= CLB_3_3_IN_pin_6_driver_mux_fanins(CLB_3_3_IN_pin_6_driver_mux_selector);
	CLB_3_3_IN_pin_7 <= CLB_3_3_IN_pin_7_driver_mux_fanins(CLB_3_3_IN_pin_7_driver_mux_selector);
	CLB_3_3_IN_pin_8 <= CLB_3_3_IN_pin_8_driver_mux_fanins(CLB_3_3_IN_pin_8_driver_mux_selector);
	CLB_3_3_IN_pin_9 <= CLB_3_3_IN_pin_9_driver_mux_fanins(CLB_3_3_IN_pin_9_driver_mux_selector);
	CLB_3_4_IN_pin_0 <= CLB_3_4_IN_pin_0_driver_mux_fanins(CLB_3_4_IN_pin_0_driver_mux_selector);
	CLB_3_4_IN_pin_1 <= CLB_3_4_IN_pin_1_driver_mux_fanins(CLB_3_4_IN_pin_1_driver_mux_selector);
	CLB_3_4_IN_pin_2 <= CLB_3_4_IN_pin_2_driver_mux_fanins(CLB_3_4_IN_pin_2_driver_mux_selector);
	CLB_3_4_IN_pin_3 <= CLB_3_4_IN_pin_3_driver_mux_fanins(CLB_3_4_IN_pin_3_driver_mux_selector);
	CLB_3_4_IN_pin_4 <= CLB_3_4_IN_pin_4_driver_mux_fanins(CLB_3_4_IN_pin_4_driver_mux_selector);
	CLB_3_4_IN_pin_5 <= CLB_3_4_IN_pin_5_driver_mux_fanins(CLB_3_4_IN_pin_5_driver_mux_selector);
	CLB_3_4_IN_pin_6 <= CLB_3_4_IN_pin_6_driver_mux_fanins(CLB_3_4_IN_pin_6_driver_mux_selector);
	CLB_3_4_IN_pin_7 <= CLB_3_4_IN_pin_7_driver_mux_fanins(CLB_3_4_IN_pin_7_driver_mux_selector);
	CLB_3_4_IN_pin_8 <= CLB_3_4_IN_pin_8_driver_mux_fanins(CLB_3_4_IN_pin_8_driver_mux_selector);
	CLB_3_4_IN_pin_9 <= CLB_3_4_IN_pin_9_driver_mux_fanins(CLB_3_4_IN_pin_9_driver_mux_selector);
	CLB_3_5_IN_pin_0 <= CLB_3_5_IN_pin_0_driver_mux_fanins(CLB_3_5_IN_pin_0_driver_mux_selector);
	CLB_3_5_IN_pin_1 <= CLB_3_5_IN_pin_1_driver_mux_fanins(CLB_3_5_IN_pin_1_driver_mux_selector);
	CLB_3_5_IN_pin_2 <= CLB_3_5_IN_pin_2_driver_mux_fanins(CLB_3_5_IN_pin_2_driver_mux_selector);
	CLB_3_5_IN_pin_3 <= CLB_3_5_IN_pin_3_driver_mux_fanins(CLB_3_5_IN_pin_3_driver_mux_selector);
	CLB_3_5_IN_pin_4 <= CLB_3_5_IN_pin_4_driver_mux_fanins(CLB_3_5_IN_pin_4_driver_mux_selector);
	CLB_3_5_IN_pin_5 <= CLB_3_5_IN_pin_5_driver_mux_fanins(CLB_3_5_IN_pin_5_driver_mux_selector);
	CLB_3_5_IN_pin_6 <= CLB_3_5_IN_pin_6_driver_mux_fanins(CLB_3_5_IN_pin_6_driver_mux_selector);
	CLB_3_5_IN_pin_7 <= CLB_3_5_IN_pin_7_driver_mux_fanins(CLB_3_5_IN_pin_7_driver_mux_selector);
	CLB_3_5_IN_pin_8 <= CLB_3_5_IN_pin_8_driver_mux_fanins(CLB_3_5_IN_pin_8_driver_mux_selector);
	CLB_3_5_IN_pin_9 <= CLB_3_5_IN_pin_9_driver_mux_fanins(CLB_3_5_IN_pin_9_driver_mux_selector);
	CLB_3_6_IN_pin_0 <= CLB_3_6_IN_pin_0_driver_mux_fanins(CLB_3_6_IN_pin_0_driver_mux_selector);
	CLB_3_6_IN_pin_1 <= CLB_3_6_IN_pin_1_driver_mux_fanins(CLB_3_6_IN_pin_1_driver_mux_selector);
	CLB_3_6_IN_pin_2 <= CLB_3_6_IN_pin_2_driver_mux_fanins(CLB_3_6_IN_pin_2_driver_mux_selector);
	CLB_3_6_IN_pin_3 <= CLB_3_6_IN_pin_3_driver_mux_fanins(CLB_3_6_IN_pin_3_driver_mux_selector);
	CLB_3_6_IN_pin_4 <= CLB_3_6_IN_pin_4_driver_mux_fanins(CLB_3_6_IN_pin_4_driver_mux_selector);
	CLB_3_6_IN_pin_5 <= CLB_3_6_IN_pin_5_driver_mux_fanins(CLB_3_6_IN_pin_5_driver_mux_selector);
	CLB_3_6_IN_pin_6 <= CLB_3_6_IN_pin_6_driver_mux_fanins(CLB_3_6_IN_pin_6_driver_mux_selector);
	CLB_3_6_IN_pin_7 <= CLB_3_6_IN_pin_7_driver_mux_fanins(CLB_3_6_IN_pin_7_driver_mux_selector);
	CLB_3_6_IN_pin_8 <= CLB_3_6_IN_pin_8_driver_mux_fanins(CLB_3_6_IN_pin_8_driver_mux_selector);
	CLB_3_6_IN_pin_9 <= CLB_3_6_IN_pin_9_driver_mux_fanins(CLB_3_6_IN_pin_9_driver_mux_selector);
	CLB_4_1_IN_pin_0 <= CLB_4_1_IN_pin_0_driver_mux_fanins(CLB_4_1_IN_pin_0_driver_mux_selector);
	CLB_4_1_IN_pin_1 <= CLB_4_1_IN_pin_1_driver_mux_fanins(CLB_4_1_IN_pin_1_driver_mux_selector);
	CLB_4_1_IN_pin_2 <= CLB_4_1_IN_pin_2_driver_mux_fanins(CLB_4_1_IN_pin_2_driver_mux_selector);
	CLB_4_1_IN_pin_3 <= CLB_4_1_IN_pin_3_driver_mux_fanins(CLB_4_1_IN_pin_3_driver_mux_selector);
	CLB_4_1_IN_pin_4 <= CLB_4_1_IN_pin_4_driver_mux_fanins(CLB_4_1_IN_pin_4_driver_mux_selector);
	CLB_4_1_IN_pin_5 <= CLB_4_1_IN_pin_5_driver_mux_fanins(CLB_4_1_IN_pin_5_driver_mux_selector);
	CLB_4_1_IN_pin_6 <= CLB_4_1_IN_pin_6_driver_mux_fanins(CLB_4_1_IN_pin_6_driver_mux_selector);
	CLB_4_1_IN_pin_7 <= CLB_4_1_IN_pin_7_driver_mux_fanins(CLB_4_1_IN_pin_7_driver_mux_selector);
	CLB_4_1_IN_pin_8 <= CLB_4_1_IN_pin_8_driver_mux_fanins(CLB_4_1_IN_pin_8_driver_mux_selector);
	CLB_4_1_IN_pin_9 <= CLB_4_1_IN_pin_9_driver_mux_fanins(CLB_4_1_IN_pin_9_driver_mux_selector);
	CLB_4_2_IN_pin_0 <= CLB_4_2_IN_pin_0_driver_mux_fanins(CLB_4_2_IN_pin_0_driver_mux_selector);
	CLB_4_2_IN_pin_1 <= CLB_4_2_IN_pin_1_driver_mux_fanins(CLB_4_2_IN_pin_1_driver_mux_selector);
	CLB_4_2_IN_pin_2 <= CLB_4_2_IN_pin_2_driver_mux_fanins(CLB_4_2_IN_pin_2_driver_mux_selector);
	CLB_4_2_IN_pin_3 <= CLB_4_2_IN_pin_3_driver_mux_fanins(CLB_4_2_IN_pin_3_driver_mux_selector);
	CLB_4_2_IN_pin_4 <= CLB_4_2_IN_pin_4_driver_mux_fanins(CLB_4_2_IN_pin_4_driver_mux_selector);
	CLB_4_2_IN_pin_5 <= CLB_4_2_IN_pin_5_driver_mux_fanins(CLB_4_2_IN_pin_5_driver_mux_selector);
	CLB_4_2_IN_pin_6 <= CLB_4_2_IN_pin_6_driver_mux_fanins(CLB_4_2_IN_pin_6_driver_mux_selector);
	CLB_4_2_IN_pin_7 <= CLB_4_2_IN_pin_7_driver_mux_fanins(CLB_4_2_IN_pin_7_driver_mux_selector);
	CLB_4_2_IN_pin_8 <= CLB_4_2_IN_pin_8_driver_mux_fanins(CLB_4_2_IN_pin_8_driver_mux_selector);
	CLB_4_2_IN_pin_9 <= CLB_4_2_IN_pin_9_driver_mux_fanins(CLB_4_2_IN_pin_9_driver_mux_selector);
	CLB_4_3_IN_pin_0 <= CLB_4_3_IN_pin_0_driver_mux_fanins(CLB_4_3_IN_pin_0_driver_mux_selector);
	CLB_4_3_IN_pin_1 <= CLB_4_3_IN_pin_1_driver_mux_fanins(CLB_4_3_IN_pin_1_driver_mux_selector);
	CLB_4_3_IN_pin_2 <= CLB_4_3_IN_pin_2_driver_mux_fanins(CLB_4_3_IN_pin_2_driver_mux_selector);
	CLB_4_3_IN_pin_3 <= CLB_4_3_IN_pin_3_driver_mux_fanins(CLB_4_3_IN_pin_3_driver_mux_selector);
	CLB_4_3_IN_pin_4 <= CLB_4_3_IN_pin_4_driver_mux_fanins(CLB_4_3_IN_pin_4_driver_mux_selector);
	CLB_4_3_IN_pin_5 <= CLB_4_3_IN_pin_5_driver_mux_fanins(CLB_4_3_IN_pin_5_driver_mux_selector);
	CLB_4_3_IN_pin_6 <= CLB_4_3_IN_pin_6_driver_mux_fanins(CLB_4_3_IN_pin_6_driver_mux_selector);
	CLB_4_3_IN_pin_7 <= CLB_4_3_IN_pin_7_driver_mux_fanins(CLB_4_3_IN_pin_7_driver_mux_selector);
	CLB_4_3_IN_pin_8 <= CLB_4_3_IN_pin_8_driver_mux_fanins(CLB_4_3_IN_pin_8_driver_mux_selector);
	CLB_4_3_IN_pin_9 <= CLB_4_3_IN_pin_9_driver_mux_fanins(CLB_4_3_IN_pin_9_driver_mux_selector);
	CLB_4_4_IN_pin_0 <= CLB_4_4_IN_pin_0_driver_mux_fanins(CLB_4_4_IN_pin_0_driver_mux_selector);
	CLB_4_4_IN_pin_1 <= CLB_4_4_IN_pin_1_driver_mux_fanins(CLB_4_4_IN_pin_1_driver_mux_selector);
	CLB_4_4_IN_pin_2 <= CLB_4_4_IN_pin_2_driver_mux_fanins(CLB_4_4_IN_pin_2_driver_mux_selector);
	CLB_4_4_IN_pin_3 <= CLB_4_4_IN_pin_3_driver_mux_fanins(CLB_4_4_IN_pin_3_driver_mux_selector);
	CLB_4_4_IN_pin_4 <= CLB_4_4_IN_pin_4_driver_mux_fanins(CLB_4_4_IN_pin_4_driver_mux_selector);
	CLB_4_4_IN_pin_5 <= CLB_4_4_IN_pin_5_driver_mux_fanins(CLB_4_4_IN_pin_5_driver_mux_selector);
	CLB_4_4_IN_pin_6 <= CLB_4_4_IN_pin_6_driver_mux_fanins(CLB_4_4_IN_pin_6_driver_mux_selector);
	CLB_4_4_IN_pin_7 <= CLB_4_4_IN_pin_7_driver_mux_fanins(CLB_4_4_IN_pin_7_driver_mux_selector);
	CLB_4_4_IN_pin_8 <= CLB_4_4_IN_pin_8_driver_mux_fanins(CLB_4_4_IN_pin_8_driver_mux_selector);
	CLB_4_4_IN_pin_9 <= CLB_4_4_IN_pin_9_driver_mux_fanins(CLB_4_4_IN_pin_9_driver_mux_selector);
	CLB_4_5_IN_pin_0 <= CLB_4_5_IN_pin_0_driver_mux_fanins(CLB_4_5_IN_pin_0_driver_mux_selector);
	CLB_4_5_IN_pin_1 <= CLB_4_5_IN_pin_1_driver_mux_fanins(CLB_4_5_IN_pin_1_driver_mux_selector);
	CLB_4_5_IN_pin_2 <= CLB_4_5_IN_pin_2_driver_mux_fanins(CLB_4_5_IN_pin_2_driver_mux_selector);
	CLB_4_5_IN_pin_3 <= CLB_4_5_IN_pin_3_driver_mux_fanins(CLB_4_5_IN_pin_3_driver_mux_selector);
	CLB_4_5_IN_pin_4 <= CLB_4_5_IN_pin_4_driver_mux_fanins(CLB_4_5_IN_pin_4_driver_mux_selector);
	CLB_4_5_IN_pin_5 <= CLB_4_5_IN_pin_5_driver_mux_fanins(CLB_4_5_IN_pin_5_driver_mux_selector);
	CLB_4_5_IN_pin_6 <= CLB_4_5_IN_pin_6_driver_mux_fanins(CLB_4_5_IN_pin_6_driver_mux_selector);
	CLB_4_5_IN_pin_7 <= CLB_4_5_IN_pin_7_driver_mux_fanins(CLB_4_5_IN_pin_7_driver_mux_selector);
	CLB_4_5_IN_pin_8 <= CLB_4_5_IN_pin_8_driver_mux_fanins(CLB_4_5_IN_pin_8_driver_mux_selector);
	CLB_4_5_IN_pin_9 <= CLB_4_5_IN_pin_9_driver_mux_fanins(CLB_4_5_IN_pin_9_driver_mux_selector);
	CLB_4_6_IN_pin_0 <= CLB_4_6_IN_pin_0_driver_mux_fanins(CLB_4_6_IN_pin_0_driver_mux_selector);
	CLB_4_6_IN_pin_1 <= CLB_4_6_IN_pin_1_driver_mux_fanins(CLB_4_6_IN_pin_1_driver_mux_selector);
	CLB_4_6_IN_pin_2 <= CLB_4_6_IN_pin_2_driver_mux_fanins(CLB_4_6_IN_pin_2_driver_mux_selector);
	CLB_4_6_IN_pin_3 <= CLB_4_6_IN_pin_3_driver_mux_fanins(CLB_4_6_IN_pin_3_driver_mux_selector);
	CLB_4_6_IN_pin_4 <= CLB_4_6_IN_pin_4_driver_mux_fanins(CLB_4_6_IN_pin_4_driver_mux_selector);
	CLB_4_6_IN_pin_5 <= CLB_4_6_IN_pin_5_driver_mux_fanins(CLB_4_6_IN_pin_5_driver_mux_selector);
	CLB_4_6_IN_pin_6 <= CLB_4_6_IN_pin_6_driver_mux_fanins(CLB_4_6_IN_pin_6_driver_mux_selector);
	CLB_4_6_IN_pin_7 <= CLB_4_6_IN_pin_7_driver_mux_fanins(CLB_4_6_IN_pin_7_driver_mux_selector);
	CLB_4_6_IN_pin_8 <= CLB_4_6_IN_pin_8_driver_mux_fanins(CLB_4_6_IN_pin_8_driver_mux_selector);
	CLB_4_6_IN_pin_9 <= CLB_4_6_IN_pin_9_driver_mux_fanins(CLB_4_6_IN_pin_9_driver_mux_selector);
	CLB_5_1_IN_pin_0 <= CLB_5_1_IN_pin_0_driver_mux_fanins(CLB_5_1_IN_pin_0_driver_mux_selector);
	CLB_5_1_IN_pin_1 <= CLB_5_1_IN_pin_1_driver_mux_fanins(CLB_5_1_IN_pin_1_driver_mux_selector);
	CLB_5_1_IN_pin_2 <= CLB_5_1_IN_pin_2_driver_mux_fanins(CLB_5_1_IN_pin_2_driver_mux_selector);
	CLB_5_1_IN_pin_3 <= CLB_5_1_IN_pin_3_driver_mux_fanins(CLB_5_1_IN_pin_3_driver_mux_selector);
	CLB_5_1_IN_pin_4 <= CLB_5_1_IN_pin_4_driver_mux_fanins(CLB_5_1_IN_pin_4_driver_mux_selector);
	CLB_5_1_IN_pin_5 <= CLB_5_1_IN_pin_5_driver_mux_fanins(CLB_5_1_IN_pin_5_driver_mux_selector);
	CLB_5_1_IN_pin_6 <= CLB_5_1_IN_pin_6_driver_mux_fanins(CLB_5_1_IN_pin_6_driver_mux_selector);
	CLB_5_1_IN_pin_7 <= CLB_5_1_IN_pin_7_driver_mux_fanins(CLB_5_1_IN_pin_7_driver_mux_selector);
	CLB_5_1_IN_pin_8 <= CLB_5_1_IN_pin_8_driver_mux_fanins(CLB_5_1_IN_pin_8_driver_mux_selector);
	CLB_5_1_IN_pin_9 <= CLB_5_1_IN_pin_9_driver_mux_fanins(CLB_5_1_IN_pin_9_driver_mux_selector);
	CLB_5_2_IN_pin_0 <= CLB_5_2_IN_pin_0_driver_mux_fanins(CLB_5_2_IN_pin_0_driver_mux_selector);
	CLB_5_2_IN_pin_1 <= CLB_5_2_IN_pin_1_driver_mux_fanins(CLB_5_2_IN_pin_1_driver_mux_selector);
	CLB_5_2_IN_pin_2 <= CLB_5_2_IN_pin_2_driver_mux_fanins(CLB_5_2_IN_pin_2_driver_mux_selector);
	CLB_5_2_IN_pin_3 <= CLB_5_2_IN_pin_3_driver_mux_fanins(CLB_5_2_IN_pin_3_driver_mux_selector);
	CLB_5_2_IN_pin_4 <= CLB_5_2_IN_pin_4_driver_mux_fanins(CLB_5_2_IN_pin_4_driver_mux_selector);
	CLB_5_2_IN_pin_5 <= CLB_5_2_IN_pin_5_driver_mux_fanins(CLB_5_2_IN_pin_5_driver_mux_selector);
	CLB_5_2_IN_pin_6 <= CLB_5_2_IN_pin_6_driver_mux_fanins(CLB_5_2_IN_pin_6_driver_mux_selector);
	CLB_5_2_IN_pin_7 <= CLB_5_2_IN_pin_7_driver_mux_fanins(CLB_5_2_IN_pin_7_driver_mux_selector);
	CLB_5_2_IN_pin_8 <= CLB_5_2_IN_pin_8_driver_mux_fanins(CLB_5_2_IN_pin_8_driver_mux_selector);
	CLB_5_2_IN_pin_9 <= CLB_5_2_IN_pin_9_driver_mux_fanins(CLB_5_2_IN_pin_9_driver_mux_selector);
	CLB_5_3_IN_pin_0 <= CLB_5_3_IN_pin_0_driver_mux_fanins(CLB_5_3_IN_pin_0_driver_mux_selector);
	CLB_5_3_IN_pin_1 <= CLB_5_3_IN_pin_1_driver_mux_fanins(CLB_5_3_IN_pin_1_driver_mux_selector);
	CLB_5_3_IN_pin_2 <= CLB_5_3_IN_pin_2_driver_mux_fanins(CLB_5_3_IN_pin_2_driver_mux_selector);
	CLB_5_3_IN_pin_3 <= CLB_5_3_IN_pin_3_driver_mux_fanins(CLB_5_3_IN_pin_3_driver_mux_selector);
	CLB_5_3_IN_pin_4 <= CLB_5_3_IN_pin_4_driver_mux_fanins(CLB_5_3_IN_pin_4_driver_mux_selector);
	CLB_5_3_IN_pin_5 <= CLB_5_3_IN_pin_5_driver_mux_fanins(CLB_5_3_IN_pin_5_driver_mux_selector);
	CLB_5_3_IN_pin_6 <= CLB_5_3_IN_pin_6_driver_mux_fanins(CLB_5_3_IN_pin_6_driver_mux_selector);
	CLB_5_3_IN_pin_7 <= CLB_5_3_IN_pin_7_driver_mux_fanins(CLB_5_3_IN_pin_7_driver_mux_selector);
	CLB_5_3_IN_pin_8 <= CLB_5_3_IN_pin_8_driver_mux_fanins(CLB_5_3_IN_pin_8_driver_mux_selector);
	CLB_5_3_IN_pin_9 <= CLB_5_3_IN_pin_9_driver_mux_fanins(CLB_5_3_IN_pin_9_driver_mux_selector);
	CLB_5_4_IN_pin_0 <= CLB_5_4_IN_pin_0_driver_mux_fanins(CLB_5_4_IN_pin_0_driver_mux_selector);
	CLB_5_4_IN_pin_1 <= CLB_5_4_IN_pin_1_driver_mux_fanins(CLB_5_4_IN_pin_1_driver_mux_selector);
	CLB_5_4_IN_pin_2 <= CLB_5_4_IN_pin_2_driver_mux_fanins(CLB_5_4_IN_pin_2_driver_mux_selector);
	CLB_5_4_IN_pin_3 <= CLB_5_4_IN_pin_3_driver_mux_fanins(CLB_5_4_IN_pin_3_driver_mux_selector);
	CLB_5_4_IN_pin_4 <= CLB_5_4_IN_pin_4_driver_mux_fanins(CLB_5_4_IN_pin_4_driver_mux_selector);
	CLB_5_4_IN_pin_5 <= CLB_5_4_IN_pin_5_driver_mux_fanins(CLB_5_4_IN_pin_5_driver_mux_selector);
	CLB_5_4_IN_pin_6 <= CLB_5_4_IN_pin_6_driver_mux_fanins(CLB_5_4_IN_pin_6_driver_mux_selector);
	CLB_5_4_IN_pin_7 <= CLB_5_4_IN_pin_7_driver_mux_fanins(CLB_5_4_IN_pin_7_driver_mux_selector);
	CLB_5_4_IN_pin_8 <= CLB_5_4_IN_pin_8_driver_mux_fanins(CLB_5_4_IN_pin_8_driver_mux_selector);
	CLB_5_4_IN_pin_9 <= CLB_5_4_IN_pin_9_driver_mux_fanins(CLB_5_4_IN_pin_9_driver_mux_selector);
	CLB_5_5_IN_pin_0 <= CLB_5_5_IN_pin_0_driver_mux_fanins(CLB_5_5_IN_pin_0_driver_mux_selector);
	CLB_5_5_IN_pin_1 <= CLB_5_5_IN_pin_1_driver_mux_fanins(CLB_5_5_IN_pin_1_driver_mux_selector);
	CLB_5_5_IN_pin_2 <= CLB_5_5_IN_pin_2_driver_mux_fanins(CLB_5_5_IN_pin_2_driver_mux_selector);
	CLB_5_5_IN_pin_3 <= CLB_5_5_IN_pin_3_driver_mux_fanins(CLB_5_5_IN_pin_3_driver_mux_selector);
	CLB_5_5_IN_pin_4 <= CLB_5_5_IN_pin_4_driver_mux_fanins(CLB_5_5_IN_pin_4_driver_mux_selector);
	CLB_5_5_IN_pin_5 <= CLB_5_5_IN_pin_5_driver_mux_fanins(CLB_5_5_IN_pin_5_driver_mux_selector);
	CLB_5_5_IN_pin_6 <= CLB_5_5_IN_pin_6_driver_mux_fanins(CLB_5_5_IN_pin_6_driver_mux_selector);
	CLB_5_5_IN_pin_7 <= CLB_5_5_IN_pin_7_driver_mux_fanins(CLB_5_5_IN_pin_7_driver_mux_selector);
	CLB_5_5_IN_pin_8 <= CLB_5_5_IN_pin_8_driver_mux_fanins(CLB_5_5_IN_pin_8_driver_mux_selector);
	CLB_5_5_IN_pin_9 <= CLB_5_5_IN_pin_9_driver_mux_fanins(CLB_5_5_IN_pin_9_driver_mux_selector);
	CLB_5_6_IN_pin_0 <= CLB_5_6_IN_pin_0_driver_mux_fanins(CLB_5_6_IN_pin_0_driver_mux_selector);
	CLB_5_6_IN_pin_1 <= CLB_5_6_IN_pin_1_driver_mux_fanins(CLB_5_6_IN_pin_1_driver_mux_selector);
	CLB_5_6_IN_pin_2 <= CLB_5_6_IN_pin_2_driver_mux_fanins(CLB_5_6_IN_pin_2_driver_mux_selector);
	CLB_5_6_IN_pin_3 <= CLB_5_6_IN_pin_3_driver_mux_fanins(CLB_5_6_IN_pin_3_driver_mux_selector);
	CLB_5_6_IN_pin_4 <= CLB_5_6_IN_pin_4_driver_mux_fanins(CLB_5_6_IN_pin_4_driver_mux_selector);
	CLB_5_6_IN_pin_5 <= CLB_5_6_IN_pin_5_driver_mux_fanins(CLB_5_6_IN_pin_5_driver_mux_selector);
	CLB_5_6_IN_pin_6 <= CLB_5_6_IN_pin_6_driver_mux_fanins(CLB_5_6_IN_pin_6_driver_mux_selector);
	CLB_5_6_IN_pin_7 <= CLB_5_6_IN_pin_7_driver_mux_fanins(CLB_5_6_IN_pin_7_driver_mux_selector);
	CLB_5_6_IN_pin_8 <= CLB_5_6_IN_pin_8_driver_mux_fanins(CLB_5_6_IN_pin_8_driver_mux_selector);
	CLB_5_6_IN_pin_9 <= CLB_5_6_IN_pin_9_driver_mux_fanins(CLB_5_6_IN_pin_9_driver_mux_selector);
	CLB_6_1_IN_pin_0 <= CLB_6_1_IN_pin_0_driver_mux_fanins(CLB_6_1_IN_pin_0_driver_mux_selector);
	CLB_6_1_IN_pin_1 <= CLB_6_1_IN_pin_1_driver_mux_fanins(CLB_6_1_IN_pin_1_driver_mux_selector);
	CLB_6_1_IN_pin_2 <= CLB_6_1_IN_pin_2_driver_mux_fanins(CLB_6_1_IN_pin_2_driver_mux_selector);
	CLB_6_1_IN_pin_3 <= CLB_6_1_IN_pin_3_driver_mux_fanins(CLB_6_1_IN_pin_3_driver_mux_selector);
	CLB_6_1_IN_pin_4 <= CLB_6_1_IN_pin_4_driver_mux_fanins(CLB_6_1_IN_pin_4_driver_mux_selector);
	CLB_6_1_IN_pin_5 <= CLB_6_1_IN_pin_5_driver_mux_fanins(CLB_6_1_IN_pin_5_driver_mux_selector);
	CLB_6_1_IN_pin_6 <= CLB_6_1_IN_pin_6_driver_mux_fanins(CLB_6_1_IN_pin_6_driver_mux_selector);
	CLB_6_1_IN_pin_7 <= CLB_6_1_IN_pin_7_driver_mux_fanins(CLB_6_1_IN_pin_7_driver_mux_selector);
	CLB_6_1_IN_pin_8 <= CLB_6_1_IN_pin_8_driver_mux_fanins(CLB_6_1_IN_pin_8_driver_mux_selector);
	CLB_6_1_IN_pin_9 <= CLB_6_1_IN_pin_9_driver_mux_fanins(CLB_6_1_IN_pin_9_driver_mux_selector);
	CLB_6_2_IN_pin_0 <= CLB_6_2_IN_pin_0_driver_mux_fanins(CLB_6_2_IN_pin_0_driver_mux_selector);
	CLB_6_2_IN_pin_1 <= CLB_6_2_IN_pin_1_driver_mux_fanins(CLB_6_2_IN_pin_1_driver_mux_selector);
	CLB_6_2_IN_pin_2 <= CLB_6_2_IN_pin_2_driver_mux_fanins(CLB_6_2_IN_pin_2_driver_mux_selector);
	CLB_6_2_IN_pin_3 <= CLB_6_2_IN_pin_3_driver_mux_fanins(CLB_6_2_IN_pin_3_driver_mux_selector);
	CLB_6_2_IN_pin_4 <= CLB_6_2_IN_pin_4_driver_mux_fanins(CLB_6_2_IN_pin_4_driver_mux_selector);
	CLB_6_2_IN_pin_5 <= CLB_6_2_IN_pin_5_driver_mux_fanins(CLB_6_2_IN_pin_5_driver_mux_selector);
	CLB_6_2_IN_pin_6 <= CLB_6_2_IN_pin_6_driver_mux_fanins(CLB_6_2_IN_pin_6_driver_mux_selector);
	CLB_6_2_IN_pin_7 <= CLB_6_2_IN_pin_7_driver_mux_fanins(CLB_6_2_IN_pin_7_driver_mux_selector);
	CLB_6_2_IN_pin_8 <= CLB_6_2_IN_pin_8_driver_mux_fanins(CLB_6_2_IN_pin_8_driver_mux_selector);
	CLB_6_2_IN_pin_9 <= CLB_6_2_IN_pin_9_driver_mux_fanins(CLB_6_2_IN_pin_9_driver_mux_selector);
	CLB_6_3_IN_pin_0 <= CLB_6_3_IN_pin_0_driver_mux_fanins(CLB_6_3_IN_pin_0_driver_mux_selector);
	CLB_6_3_IN_pin_1 <= CLB_6_3_IN_pin_1_driver_mux_fanins(CLB_6_3_IN_pin_1_driver_mux_selector);
	CLB_6_3_IN_pin_2 <= CLB_6_3_IN_pin_2_driver_mux_fanins(CLB_6_3_IN_pin_2_driver_mux_selector);
	CLB_6_3_IN_pin_3 <= CLB_6_3_IN_pin_3_driver_mux_fanins(CLB_6_3_IN_pin_3_driver_mux_selector);
	CLB_6_3_IN_pin_4 <= CLB_6_3_IN_pin_4_driver_mux_fanins(CLB_6_3_IN_pin_4_driver_mux_selector);
	CLB_6_3_IN_pin_5 <= CLB_6_3_IN_pin_5_driver_mux_fanins(CLB_6_3_IN_pin_5_driver_mux_selector);
	CLB_6_3_IN_pin_6 <= CLB_6_3_IN_pin_6_driver_mux_fanins(CLB_6_3_IN_pin_6_driver_mux_selector);
	CLB_6_3_IN_pin_7 <= CLB_6_3_IN_pin_7_driver_mux_fanins(CLB_6_3_IN_pin_7_driver_mux_selector);
	CLB_6_3_IN_pin_8 <= CLB_6_3_IN_pin_8_driver_mux_fanins(CLB_6_3_IN_pin_8_driver_mux_selector);
	CLB_6_3_IN_pin_9 <= CLB_6_3_IN_pin_9_driver_mux_fanins(CLB_6_3_IN_pin_9_driver_mux_selector);
	CLB_6_4_IN_pin_0 <= CLB_6_4_IN_pin_0_driver_mux_fanins(CLB_6_4_IN_pin_0_driver_mux_selector);
	CLB_6_4_IN_pin_1 <= CLB_6_4_IN_pin_1_driver_mux_fanins(CLB_6_4_IN_pin_1_driver_mux_selector);
	CLB_6_4_IN_pin_2 <= CLB_6_4_IN_pin_2_driver_mux_fanins(CLB_6_4_IN_pin_2_driver_mux_selector);
	CLB_6_4_IN_pin_3 <= CLB_6_4_IN_pin_3_driver_mux_fanins(CLB_6_4_IN_pin_3_driver_mux_selector);
	CLB_6_4_IN_pin_4 <= CLB_6_4_IN_pin_4_driver_mux_fanins(CLB_6_4_IN_pin_4_driver_mux_selector);
	CLB_6_4_IN_pin_5 <= CLB_6_4_IN_pin_5_driver_mux_fanins(CLB_6_4_IN_pin_5_driver_mux_selector);
	CLB_6_4_IN_pin_6 <= CLB_6_4_IN_pin_6_driver_mux_fanins(CLB_6_4_IN_pin_6_driver_mux_selector);
	CLB_6_4_IN_pin_7 <= CLB_6_4_IN_pin_7_driver_mux_fanins(CLB_6_4_IN_pin_7_driver_mux_selector);
	CLB_6_4_IN_pin_8 <= CLB_6_4_IN_pin_8_driver_mux_fanins(CLB_6_4_IN_pin_8_driver_mux_selector);
	CLB_6_4_IN_pin_9 <= CLB_6_4_IN_pin_9_driver_mux_fanins(CLB_6_4_IN_pin_9_driver_mux_selector);
	CLB_6_5_IN_pin_0 <= CLB_6_5_IN_pin_0_driver_mux_fanins(CLB_6_5_IN_pin_0_driver_mux_selector);
	CLB_6_5_IN_pin_1 <= CLB_6_5_IN_pin_1_driver_mux_fanins(CLB_6_5_IN_pin_1_driver_mux_selector);
	CLB_6_5_IN_pin_2 <= CLB_6_5_IN_pin_2_driver_mux_fanins(CLB_6_5_IN_pin_2_driver_mux_selector);
	CLB_6_5_IN_pin_3 <= CLB_6_5_IN_pin_3_driver_mux_fanins(CLB_6_5_IN_pin_3_driver_mux_selector);
	CLB_6_5_IN_pin_4 <= CLB_6_5_IN_pin_4_driver_mux_fanins(CLB_6_5_IN_pin_4_driver_mux_selector);
	CLB_6_5_IN_pin_5 <= CLB_6_5_IN_pin_5_driver_mux_fanins(CLB_6_5_IN_pin_5_driver_mux_selector);
	CLB_6_5_IN_pin_6 <= CLB_6_5_IN_pin_6_driver_mux_fanins(CLB_6_5_IN_pin_6_driver_mux_selector);
	CLB_6_5_IN_pin_7 <= CLB_6_5_IN_pin_7_driver_mux_fanins(CLB_6_5_IN_pin_7_driver_mux_selector);
	CLB_6_5_IN_pin_8 <= CLB_6_5_IN_pin_8_driver_mux_fanins(CLB_6_5_IN_pin_8_driver_mux_selector);
	CLB_6_5_IN_pin_9 <= CLB_6_5_IN_pin_9_driver_mux_fanins(CLB_6_5_IN_pin_9_driver_mux_selector);
	CLB_6_6_IN_pin_0 <= CLB_6_6_IN_pin_0_driver_mux_fanins(CLB_6_6_IN_pin_0_driver_mux_selector);
	CLB_6_6_IN_pin_1 <= CLB_6_6_IN_pin_1_driver_mux_fanins(CLB_6_6_IN_pin_1_driver_mux_selector);
	CLB_6_6_IN_pin_2 <= CLB_6_6_IN_pin_2_driver_mux_fanins(CLB_6_6_IN_pin_2_driver_mux_selector);
	CLB_6_6_IN_pin_3 <= CLB_6_6_IN_pin_3_driver_mux_fanins(CLB_6_6_IN_pin_3_driver_mux_selector);
	CLB_6_6_IN_pin_4 <= CLB_6_6_IN_pin_4_driver_mux_fanins(CLB_6_6_IN_pin_4_driver_mux_selector);
	CLB_6_6_IN_pin_5 <= CLB_6_6_IN_pin_5_driver_mux_fanins(CLB_6_6_IN_pin_5_driver_mux_selector);
	CLB_6_6_IN_pin_6 <= CLB_6_6_IN_pin_6_driver_mux_fanins(CLB_6_6_IN_pin_6_driver_mux_selector);
	CLB_6_6_IN_pin_7 <= CLB_6_6_IN_pin_7_driver_mux_fanins(CLB_6_6_IN_pin_7_driver_mux_selector);
	CLB_6_6_IN_pin_8 <= CLB_6_6_IN_pin_8_driver_mux_fanins(CLB_6_6_IN_pin_8_driver_mux_selector);
	CLB_6_6_IN_pin_9 <= CLB_6_6_IN_pin_9_driver_mux_fanins(CLB_6_6_IN_pin_9_driver_mux_selector);
	CLB_7_1_IN_pin_0 <= CLB_7_1_IN_pin_0_driver_mux_fanins(CLB_7_1_IN_pin_0_driver_mux_selector);
	CLB_7_1_IN_pin_1 <= CLB_7_1_IN_pin_1_driver_mux_fanins(CLB_7_1_IN_pin_1_driver_mux_selector);
	CLB_7_1_IN_pin_2 <= CLB_7_1_IN_pin_2_driver_mux_fanins(CLB_7_1_IN_pin_2_driver_mux_selector);
	CLB_7_1_IN_pin_3 <= CLB_7_1_IN_pin_3_driver_mux_fanins(CLB_7_1_IN_pin_3_driver_mux_selector);
	CLB_7_1_IN_pin_4 <= CLB_7_1_IN_pin_4_driver_mux_fanins(CLB_7_1_IN_pin_4_driver_mux_selector);
	CLB_7_1_IN_pin_5 <= CLB_7_1_IN_pin_5_driver_mux_fanins(CLB_7_1_IN_pin_5_driver_mux_selector);
	CLB_7_1_IN_pin_6 <= CLB_7_1_IN_pin_6_driver_mux_fanins(CLB_7_1_IN_pin_6_driver_mux_selector);
	CLB_7_1_IN_pin_7 <= CLB_7_1_IN_pin_7_driver_mux_fanins(CLB_7_1_IN_pin_7_driver_mux_selector);
	CLB_7_1_IN_pin_8 <= CLB_7_1_IN_pin_8_driver_mux_fanins(CLB_7_1_IN_pin_8_driver_mux_selector);
	CLB_7_1_IN_pin_9 <= CLB_7_1_IN_pin_9_driver_mux_fanins(CLB_7_1_IN_pin_9_driver_mux_selector);
	CLB_7_2_IN_pin_0 <= CLB_7_2_IN_pin_0_driver_mux_fanins(CLB_7_2_IN_pin_0_driver_mux_selector);
	CLB_7_2_IN_pin_1 <= CLB_7_2_IN_pin_1_driver_mux_fanins(CLB_7_2_IN_pin_1_driver_mux_selector);
	CLB_7_2_IN_pin_2 <= CLB_7_2_IN_pin_2_driver_mux_fanins(CLB_7_2_IN_pin_2_driver_mux_selector);
	CLB_7_2_IN_pin_3 <= CLB_7_2_IN_pin_3_driver_mux_fanins(CLB_7_2_IN_pin_3_driver_mux_selector);
	CLB_7_2_IN_pin_4 <= CLB_7_2_IN_pin_4_driver_mux_fanins(CLB_7_2_IN_pin_4_driver_mux_selector);
	CLB_7_2_IN_pin_5 <= CLB_7_2_IN_pin_5_driver_mux_fanins(CLB_7_2_IN_pin_5_driver_mux_selector);
	CLB_7_2_IN_pin_6 <= CLB_7_2_IN_pin_6_driver_mux_fanins(CLB_7_2_IN_pin_6_driver_mux_selector);
	CLB_7_2_IN_pin_7 <= CLB_7_2_IN_pin_7_driver_mux_fanins(CLB_7_2_IN_pin_7_driver_mux_selector);
	CLB_7_2_IN_pin_8 <= CLB_7_2_IN_pin_8_driver_mux_fanins(CLB_7_2_IN_pin_8_driver_mux_selector);
	CLB_7_2_IN_pin_9 <= CLB_7_2_IN_pin_9_driver_mux_fanins(CLB_7_2_IN_pin_9_driver_mux_selector);
	CLB_7_3_IN_pin_0 <= CLB_7_3_IN_pin_0_driver_mux_fanins(CLB_7_3_IN_pin_0_driver_mux_selector);
	CLB_7_3_IN_pin_1 <= CLB_7_3_IN_pin_1_driver_mux_fanins(CLB_7_3_IN_pin_1_driver_mux_selector);
	CLB_7_3_IN_pin_2 <= CLB_7_3_IN_pin_2_driver_mux_fanins(CLB_7_3_IN_pin_2_driver_mux_selector);
	CLB_7_3_IN_pin_3 <= CLB_7_3_IN_pin_3_driver_mux_fanins(CLB_7_3_IN_pin_3_driver_mux_selector);
	CLB_7_3_IN_pin_4 <= CLB_7_3_IN_pin_4_driver_mux_fanins(CLB_7_3_IN_pin_4_driver_mux_selector);
	CLB_7_3_IN_pin_5 <= CLB_7_3_IN_pin_5_driver_mux_fanins(CLB_7_3_IN_pin_5_driver_mux_selector);
	CLB_7_3_IN_pin_6 <= CLB_7_3_IN_pin_6_driver_mux_fanins(CLB_7_3_IN_pin_6_driver_mux_selector);
	CLB_7_3_IN_pin_7 <= CLB_7_3_IN_pin_7_driver_mux_fanins(CLB_7_3_IN_pin_7_driver_mux_selector);
	CLB_7_3_IN_pin_8 <= CLB_7_3_IN_pin_8_driver_mux_fanins(CLB_7_3_IN_pin_8_driver_mux_selector);
	CLB_7_3_IN_pin_9 <= CLB_7_3_IN_pin_9_driver_mux_fanins(CLB_7_3_IN_pin_9_driver_mux_selector);
	CLB_7_4_IN_pin_0 <= CLB_7_4_IN_pin_0_driver_mux_fanins(CLB_7_4_IN_pin_0_driver_mux_selector);
	CLB_7_4_IN_pin_1 <= CLB_7_4_IN_pin_1_driver_mux_fanins(CLB_7_4_IN_pin_1_driver_mux_selector);
	CLB_7_4_IN_pin_2 <= CLB_7_4_IN_pin_2_driver_mux_fanins(CLB_7_4_IN_pin_2_driver_mux_selector);
	CLB_7_4_IN_pin_3 <= CLB_7_4_IN_pin_3_driver_mux_fanins(CLB_7_4_IN_pin_3_driver_mux_selector);
	CLB_7_4_IN_pin_4 <= CLB_7_4_IN_pin_4_driver_mux_fanins(CLB_7_4_IN_pin_4_driver_mux_selector);
	CLB_7_4_IN_pin_5 <= CLB_7_4_IN_pin_5_driver_mux_fanins(CLB_7_4_IN_pin_5_driver_mux_selector);
	CLB_7_4_IN_pin_6 <= CLB_7_4_IN_pin_6_driver_mux_fanins(CLB_7_4_IN_pin_6_driver_mux_selector);
	CLB_7_4_IN_pin_7 <= CLB_7_4_IN_pin_7_driver_mux_fanins(CLB_7_4_IN_pin_7_driver_mux_selector);
	CLB_7_4_IN_pin_8 <= CLB_7_4_IN_pin_8_driver_mux_fanins(CLB_7_4_IN_pin_8_driver_mux_selector);
	CLB_7_4_IN_pin_9 <= CLB_7_4_IN_pin_9_driver_mux_fanins(CLB_7_4_IN_pin_9_driver_mux_selector);
	CLB_7_5_IN_pin_0 <= CLB_7_5_IN_pin_0_driver_mux_fanins(CLB_7_5_IN_pin_0_driver_mux_selector);
	CLB_7_5_IN_pin_1 <= CLB_7_5_IN_pin_1_driver_mux_fanins(CLB_7_5_IN_pin_1_driver_mux_selector);
	CLB_7_5_IN_pin_2 <= CLB_7_5_IN_pin_2_driver_mux_fanins(CLB_7_5_IN_pin_2_driver_mux_selector);
	CLB_7_5_IN_pin_3 <= CLB_7_5_IN_pin_3_driver_mux_fanins(CLB_7_5_IN_pin_3_driver_mux_selector);
	CLB_7_5_IN_pin_4 <= CLB_7_5_IN_pin_4_driver_mux_fanins(CLB_7_5_IN_pin_4_driver_mux_selector);
	CLB_7_5_IN_pin_5 <= CLB_7_5_IN_pin_5_driver_mux_fanins(CLB_7_5_IN_pin_5_driver_mux_selector);
	CLB_7_5_IN_pin_6 <= CLB_7_5_IN_pin_6_driver_mux_fanins(CLB_7_5_IN_pin_6_driver_mux_selector);
	CLB_7_5_IN_pin_7 <= CLB_7_5_IN_pin_7_driver_mux_fanins(CLB_7_5_IN_pin_7_driver_mux_selector);
	CLB_7_5_IN_pin_8 <= CLB_7_5_IN_pin_8_driver_mux_fanins(CLB_7_5_IN_pin_8_driver_mux_selector);
	CLB_7_5_IN_pin_9 <= CLB_7_5_IN_pin_9_driver_mux_fanins(CLB_7_5_IN_pin_9_driver_mux_selector);
	CLB_7_6_IN_pin_0 <= CLB_7_6_IN_pin_0_driver_mux_fanins(CLB_7_6_IN_pin_0_driver_mux_selector);
	CLB_7_6_IN_pin_1 <= CLB_7_6_IN_pin_1_driver_mux_fanins(CLB_7_6_IN_pin_1_driver_mux_selector);
	CLB_7_6_IN_pin_2 <= CLB_7_6_IN_pin_2_driver_mux_fanins(CLB_7_6_IN_pin_2_driver_mux_selector);
	CLB_7_6_IN_pin_3 <= CLB_7_6_IN_pin_3_driver_mux_fanins(CLB_7_6_IN_pin_3_driver_mux_selector);
	CLB_7_6_IN_pin_4 <= CLB_7_6_IN_pin_4_driver_mux_fanins(CLB_7_6_IN_pin_4_driver_mux_selector);
	CLB_7_6_IN_pin_5 <= CLB_7_6_IN_pin_5_driver_mux_fanins(CLB_7_6_IN_pin_5_driver_mux_selector);
	CLB_7_6_IN_pin_6 <= CLB_7_6_IN_pin_6_driver_mux_fanins(CLB_7_6_IN_pin_6_driver_mux_selector);
	CLB_7_6_IN_pin_7 <= CLB_7_6_IN_pin_7_driver_mux_fanins(CLB_7_6_IN_pin_7_driver_mux_selector);
	CLB_7_6_IN_pin_8 <= CLB_7_6_IN_pin_8_driver_mux_fanins(CLB_7_6_IN_pin_8_driver_mux_selector);
	CLB_7_6_IN_pin_9 <= CLB_7_6_IN_pin_9_driver_mux_fanins(CLB_7_6_IN_pin_9_driver_mux_selector);
	CLB_8_1_IN_pin_0 <= CLB_8_1_IN_pin_0_driver_mux_fanins(CLB_8_1_IN_pin_0_driver_mux_selector);
	CLB_8_1_IN_pin_1 <= CLB_8_1_IN_pin_1_driver_mux_fanins(CLB_8_1_IN_pin_1_driver_mux_selector);
	CLB_8_1_IN_pin_2 <= CLB_8_1_IN_pin_2_driver_mux_fanins(CLB_8_1_IN_pin_2_driver_mux_selector);
	CLB_8_1_IN_pin_3 <= CLB_8_1_IN_pin_3_driver_mux_fanins(CLB_8_1_IN_pin_3_driver_mux_selector);
	CLB_8_1_IN_pin_4 <= CLB_8_1_IN_pin_4_driver_mux_fanins(CLB_8_1_IN_pin_4_driver_mux_selector);
	CLB_8_1_IN_pin_5 <= CLB_8_1_IN_pin_5_driver_mux_fanins(CLB_8_1_IN_pin_5_driver_mux_selector);
	CLB_8_1_IN_pin_6 <= CLB_8_1_IN_pin_6_driver_mux_fanins(CLB_8_1_IN_pin_6_driver_mux_selector);
	CLB_8_1_IN_pin_7 <= CLB_8_1_IN_pin_7_driver_mux_fanins(CLB_8_1_IN_pin_7_driver_mux_selector);
	CLB_8_1_IN_pin_8 <= CLB_8_1_IN_pin_8_driver_mux_fanins(CLB_8_1_IN_pin_8_driver_mux_selector);
	CLB_8_1_IN_pin_9 <= CLB_8_1_IN_pin_9_driver_mux_fanins(CLB_8_1_IN_pin_9_driver_mux_selector);
	CLB_8_2_IN_pin_0 <= CLB_8_2_IN_pin_0_driver_mux_fanins(CLB_8_2_IN_pin_0_driver_mux_selector);
	CLB_8_2_IN_pin_1 <= CLB_8_2_IN_pin_1_driver_mux_fanins(CLB_8_2_IN_pin_1_driver_mux_selector);
	CLB_8_2_IN_pin_2 <= CLB_8_2_IN_pin_2_driver_mux_fanins(CLB_8_2_IN_pin_2_driver_mux_selector);
	CLB_8_2_IN_pin_3 <= CLB_8_2_IN_pin_3_driver_mux_fanins(CLB_8_2_IN_pin_3_driver_mux_selector);
	CLB_8_2_IN_pin_4 <= CLB_8_2_IN_pin_4_driver_mux_fanins(CLB_8_2_IN_pin_4_driver_mux_selector);
	CLB_8_2_IN_pin_5 <= CLB_8_2_IN_pin_5_driver_mux_fanins(CLB_8_2_IN_pin_5_driver_mux_selector);
	CLB_8_2_IN_pin_6 <= CLB_8_2_IN_pin_6_driver_mux_fanins(CLB_8_2_IN_pin_6_driver_mux_selector);
	CLB_8_2_IN_pin_7 <= CLB_8_2_IN_pin_7_driver_mux_fanins(CLB_8_2_IN_pin_7_driver_mux_selector);
	CLB_8_2_IN_pin_8 <= CLB_8_2_IN_pin_8_driver_mux_fanins(CLB_8_2_IN_pin_8_driver_mux_selector);
	CLB_8_2_IN_pin_9 <= CLB_8_2_IN_pin_9_driver_mux_fanins(CLB_8_2_IN_pin_9_driver_mux_selector);
	CLB_8_3_IN_pin_0 <= CLB_8_3_IN_pin_0_driver_mux_fanins(CLB_8_3_IN_pin_0_driver_mux_selector);
	CLB_8_3_IN_pin_1 <= CLB_8_3_IN_pin_1_driver_mux_fanins(CLB_8_3_IN_pin_1_driver_mux_selector);
	CLB_8_3_IN_pin_2 <= CLB_8_3_IN_pin_2_driver_mux_fanins(CLB_8_3_IN_pin_2_driver_mux_selector);
	CLB_8_3_IN_pin_3 <= CLB_8_3_IN_pin_3_driver_mux_fanins(CLB_8_3_IN_pin_3_driver_mux_selector);
	CLB_8_3_IN_pin_4 <= CLB_8_3_IN_pin_4_driver_mux_fanins(CLB_8_3_IN_pin_4_driver_mux_selector);
	CLB_8_3_IN_pin_5 <= CLB_8_3_IN_pin_5_driver_mux_fanins(CLB_8_3_IN_pin_5_driver_mux_selector);
	CLB_8_3_IN_pin_6 <= CLB_8_3_IN_pin_6_driver_mux_fanins(CLB_8_3_IN_pin_6_driver_mux_selector);
	CLB_8_3_IN_pin_7 <= CLB_8_3_IN_pin_7_driver_mux_fanins(CLB_8_3_IN_pin_7_driver_mux_selector);
	CLB_8_3_IN_pin_8 <= CLB_8_3_IN_pin_8_driver_mux_fanins(CLB_8_3_IN_pin_8_driver_mux_selector);
	CLB_8_3_IN_pin_9 <= CLB_8_3_IN_pin_9_driver_mux_fanins(CLB_8_3_IN_pin_9_driver_mux_selector);
	CLB_8_4_IN_pin_0 <= CLB_8_4_IN_pin_0_driver_mux_fanins(CLB_8_4_IN_pin_0_driver_mux_selector);
	CLB_8_4_IN_pin_1 <= CLB_8_4_IN_pin_1_driver_mux_fanins(CLB_8_4_IN_pin_1_driver_mux_selector);
	CLB_8_4_IN_pin_2 <= CLB_8_4_IN_pin_2_driver_mux_fanins(CLB_8_4_IN_pin_2_driver_mux_selector);
	CLB_8_4_IN_pin_3 <= CLB_8_4_IN_pin_3_driver_mux_fanins(CLB_8_4_IN_pin_3_driver_mux_selector);
	CLB_8_4_IN_pin_4 <= CLB_8_4_IN_pin_4_driver_mux_fanins(CLB_8_4_IN_pin_4_driver_mux_selector);
	CLB_8_4_IN_pin_5 <= CLB_8_4_IN_pin_5_driver_mux_fanins(CLB_8_4_IN_pin_5_driver_mux_selector);
	CLB_8_4_IN_pin_6 <= CLB_8_4_IN_pin_6_driver_mux_fanins(CLB_8_4_IN_pin_6_driver_mux_selector);
	CLB_8_4_IN_pin_7 <= CLB_8_4_IN_pin_7_driver_mux_fanins(CLB_8_4_IN_pin_7_driver_mux_selector);
	CLB_8_4_IN_pin_8 <= CLB_8_4_IN_pin_8_driver_mux_fanins(CLB_8_4_IN_pin_8_driver_mux_selector);
	CLB_8_4_IN_pin_9 <= CLB_8_4_IN_pin_9_driver_mux_fanins(CLB_8_4_IN_pin_9_driver_mux_selector);
	CLB_8_5_IN_pin_0 <= CLB_8_5_IN_pin_0_driver_mux_fanins(CLB_8_5_IN_pin_0_driver_mux_selector);
	CLB_8_5_IN_pin_1 <= CLB_8_5_IN_pin_1_driver_mux_fanins(CLB_8_5_IN_pin_1_driver_mux_selector);
	CLB_8_5_IN_pin_2 <= CLB_8_5_IN_pin_2_driver_mux_fanins(CLB_8_5_IN_pin_2_driver_mux_selector);
	CLB_8_5_IN_pin_3 <= CLB_8_5_IN_pin_3_driver_mux_fanins(CLB_8_5_IN_pin_3_driver_mux_selector);
	CLB_8_5_IN_pin_4 <= CLB_8_5_IN_pin_4_driver_mux_fanins(CLB_8_5_IN_pin_4_driver_mux_selector);
	CLB_8_5_IN_pin_5 <= CLB_8_5_IN_pin_5_driver_mux_fanins(CLB_8_5_IN_pin_5_driver_mux_selector);
	CLB_8_5_IN_pin_6 <= CLB_8_5_IN_pin_6_driver_mux_fanins(CLB_8_5_IN_pin_6_driver_mux_selector);
	CLB_8_5_IN_pin_7 <= CLB_8_5_IN_pin_7_driver_mux_fanins(CLB_8_5_IN_pin_7_driver_mux_selector);
	CLB_8_5_IN_pin_8 <= CLB_8_5_IN_pin_8_driver_mux_fanins(CLB_8_5_IN_pin_8_driver_mux_selector);
	CLB_8_5_IN_pin_9 <= CLB_8_5_IN_pin_9_driver_mux_fanins(CLB_8_5_IN_pin_9_driver_mux_selector);
	CLB_8_6_IN_pin_0 <= CLB_8_6_IN_pin_0_driver_mux_fanins(CLB_8_6_IN_pin_0_driver_mux_selector);
	CLB_8_6_IN_pin_1 <= CLB_8_6_IN_pin_1_driver_mux_fanins(CLB_8_6_IN_pin_1_driver_mux_selector);
	CLB_8_6_IN_pin_2 <= CLB_8_6_IN_pin_2_driver_mux_fanins(CLB_8_6_IN_pin_2_driver_mux_selector);
	CLB_8_6_IN_pin_3 <= CLB_8_6_IN_pin_3_driver_mux_fanins(CLB_8_6_IN_pin_3_driver_mux_selector);
	CLB_8_6_IN_pin_4 <= CLB_8_6_IN_pin_4_driver_mux_fanins(CLB_8_6_IN_pin_4_driver_mux_selector);
	CLB_8_6_IN_pin_5 <= CLB_8_6_IN_pin_5_driver_mux_fanins(CLB_8_6_IN_pin_5_driver_mux_selector);
	CLB_8_6_IN_pin_6 <= CLB_8_6_IN_pin_6_driver_mux_fanins(CLB_8_6_IN_pin_6_driver_mux_selector);
	CLB_8_6_IN_pin_7 <= CLB_8_6_IN_pin_7_driver_mux_fanins(CLB_8_6_IN_pin_7_driver_mux_selector);
	CLB_8_6_IN_pin_8 <= CLB_8_6_IN_pin_8_driver_mux_fanins(CLB_8_6_IN_pin_8_driver_mux_selector);
	CLB_8_6_IN_pin_9 <= CLB_8_6_IN_pin_9_driver_mux_fanins(CLB_8_6_IN_pin_9_driver_mux_selector);
	IO_0_1_IN_pin_0  <= IO_0_1_IN_pin_0_driver_mux_fanins(IO_0_1_IN_pin_0_driver_mux_selector);
	IO_0_1_IN_pin_1  <= IO_0_1_IN_pin_1_driver_mux_fanins(IO_0_1_IN_pin_1_driver_mux_selector);
	IO_0_2_IN_pin_0  <= IO_0_2_IN_pin_0_driver_mux_fanins(IO_0_2_IN_pin_0_driver_mux_selector);
	IO_0_2_IN_pin_1  <= IO_0_2_IN_pin_1_driver_mux_fanins(IO_0_2_IN_pin_1_driver_mux_selector);
	IO_0_3_IN_pin_0  <= IO_0_3_IN_pin_0_driver_mux_fanins(IO_0_3_IN_pin_0_driver_mux_selector);
	IO_0_3_IN_pin_1  <= IO_0_3_IN_pin_1_driver_mux_fanins(IO_0_3_IN_pin_1_driver_mux_selector);
	IO_0_4_IN_pin_0  <= IO_0_4_IN_pin_0_driver_mux_fanins(IO_0_4_IN_pin_0_driver_mux_selector);
	IO_0_4_IN_pin_1  <= IO_0_4_IN_pin_1_driver_mux_fanins(IO_0_4_IN_pin_1_driver_mux_selector);
	IO_0_5_IN_pin_0  <= IO_0_5_IN_pin_0_driver_mux_fanins(IO_0_5_IN_pin_0_driver_mux_selector);
	IO_0_5_IN_pin_1  <= IO_0_5_IN_pin_1_driver_mux_fanins(IO_0_5_IN_pin_1_driver_mux_selector);
	IO_0_6_IN_pin_0  <= IO_0_6_IN_pin_0_driver_mux_fanins(IO_0_6_IN_pin_0_driver_mux_selector);
	IO_0_6_IN_pin_1  <= IO_0_6_IN_pin_1_driver_mux_fanins(IO_0_6_IN_pin_1_driver_mux_selector);
	IO_1_0_IN_pin_0  <= IO_1_0_IN_pin_0_driver_mux_fanins(IO_1_0_IN_pin_0_driver_mux_selector);
	IO_1_0_IN_pin_1  <= IO_1_0_IN_pin_1_driver_mux_fanins(IO_1_0_IN_pin_1_driver_mux_selector);
	IO_1_7_IN_pin_0  <= IO_1_7_IN_pin_0_driver_mux_fanins(IO_1_7_IN_pin_0_driver_mux_selector);
	IO_1_7_IN_pin_1  <= IO_1_7_IN_pin_1_driver_mux_fanins(IO_1_7_IN_pin_1_driver_mux_selector);
	IO_2_0_IN_pin_0  <= IO_2_0_IN_pin_0_driver_mux_fanins(IO_2_0_IN_pin_0_driver_mux_selector);
	IO_2_0_IN_pin_1  <= IO_2_0_IN_pin_1_driver_mux_fanins(IO_2_0_IN_pin_1_driver_mux_selector);
	IO_2_7_IN_pin_0  <= IO_2_7_IN_pin_0_driver_mux_fanins(IO_2_7_IN_pin_0_driver_mux_selector);
	IO_2_7_IN_pin_1  <= IO_2_7_IN_pin_1_driver_mux_fanins(IO_2_7_IN_pin_1_driver_mux_selector);
	IO_3_0_IN_pin_0  <= IO_3_0_IN_pin_0_driver_mux_fanins(IO_3_0_IN_pin_0_driver_mux_selector);
	IO_3_0_IN_pin_1  <= IO_3_0_IN_pin_1_driver_mux_fanins(IO_3_0_IN_pin_1_driver_mux_selector);
	IO_3_7_IN_pin_0  <= IO_3_7_IN_pin_0_driver_mux_fanins(IO_3_7_IN_pin_0_driver_mux_selector);
	IO_3_7_IN_pin_1  <= IO_3_7_IN_pin_1_driver_mux_fanins(IO_3_7_IN_pin_1_driver_mux_selector);
	IO_4_0_IN_pin_0  <= IO_4_0_IN_pin_0_driver_mux_fanins(IO_4_0_IN_pin_0_driver_mux_selector);
	IO_4_0_IN_pin_1  <= IO_4_0_IN_pin_1_driver_mux_fanins(IO_4_0_IN_pin_1_driver_mux_selector);
	IO_4_7_IN_pin_0  <= IO_4_7_IN_pin_0_driver_mux_fanins(IO_4_7_IN_pin_0_driver_mux_selector);
	IO_4_7_IN_pin_1  <= IO_4_7_IN_pin_1_driver_mux_fanins(IO_4_7_IN_pin_1_driver_mux_selector);
	IO_5_0_IN_pin_0  <= IO_5_0_IN_pin_0_driver_mux_fanins(IO_5_0_IN_pin_0_driver_mux_selector);
	IO_5_0_IN_pin_1  <= IO_5_0_IN_pin_1_driver_mux_fanins(IO_5_0_IN_pin_1_driver_mux_selector);
	IO_5_7_IN_pin_0  <= IO_5_7_IN_pin_0_driver_mux_fanins(IO_5_7_IN_pin_0_driver_mux_selector);
	IO_5_7_IN_pin_1  <= IO_5_7_IN_pin_1_driver_mux_fanins(IO_5_7_IN_pin_1_driver_mux_selector);
	IO_6_0_IN_pin_0  <= IO_6_0_IN_pin_0_driver_mux_fanins(IO_6_0_IN_pin_0_driver_mux_selector);
	IO_6_0_IN_pin_1  <= IO_6_0_IN_pin_1_driver_mux_fanins(IO_6_0_IN_pin_1_driver_mux_selector);
	IO_6_7_IN_pin_0  <= IO_6_7_IN_pin_0_driver_mux_fanins(IO_6_7_IN_pin_0_driver_mux_selector);
	IO_6_7_IN_pin_1  <= IO_6_7_IN_pin_1_driver_mux_fanins(IO_6_7_IN_pin_1_driver_mux_selector);
	IO_7_0_IN_pin_0  <= IO_7_0_IN_pin_0_driver_mux_fanins(IO_7_0_IN_pin_0_driver_mux_selector);
	IO_7_0_IN_pin_1  <= IO_7_0_IN_pin_1_driver_mux_fanins(IO_7_0_IN_pin_1_driver_mux_selector);
	IO_7_7_IN_pin_0  <= IO_7_7_IN_pin_0_driver_mux_fanins(IO_7_7_IN_pin_0_driver_mux_selector);
	IO_7_7_IN_pin_1  <= IO_7_7_IN_pin_1_driver_mux_fanins(IO_7_7_IN_pin_1_driver_mux_selector);
	IO_8_0_IN_pin_0  <= IO_8_0_IN_pin_0_driver_mux_fanins(IO_8_0_IN_pin_0_driver_mux_selector);
	IO_8_0_IN_pin_1  <= IO_8_0_IN_pin_1_driver_mux_fanins(IO_8_0_IN_pin_1_driver_mux_selector);
	IO_8_7_IN_pin_0  <= IO_8_7_IN_pin_0_driver_mux_fanins(IO_8_7_IN_pin_0_driver_mux_selector);
	IO_8_7_IN_pin_1  <= IO_8_7_IN_pin_1_driver_mux_fanins(IO_8_7_IN_pin_1_driver_mux_selector);
	IO_9_1_IN_pin_0  <= IO_9_1_IN_pin_0_driver_mux_fanins(IO_9_1_IN_pin_0_driver_mux_selector);
	IO_9_1_IN_pin_1  <= IO_9_1_IN_pin_1_driver_mux_fanins(IO_9_1_IN_pin_1_driver_mux_selector);
	IO_9_2_IN_pin_0  <= IO_9_2_IN_pin_0_driver_mux_fanins(IO_9_2_IN_pin_0_driver_mux_selector);
	IO_9_2_IN_pin_1  <= IO_9_2_IN_pin_1_driver_mux_fanins(IO_9_2_IN_pin_1_driver_mux_selector);
	IO_9_3_IN_pin_0  <= IO_9_3_IN_pin_0_driver_mux_fanins(IO_9_3_IN_pin_0_driver_mux_selector);
	IO_9_3_IN_pin_1  <= IO_9_3_IN_pin_1_driver_mux_fanins(IO_9_3_IN_pin_1_driver_mux_selector);
	IO_9_4_IN_pin_0  <= IO_9_4_IN_pin_0_driver_mux_fanins(IO_9_4_IN_pin_0_driver_mux_selector);
	IO_9_4_IN_pin_1  <= IO_9_4_IN_pin_1_driver_mux_fanins(IO_9_4_IN_pin_1_driver_mux_selector);
	IO_9_5_IN_pin_0  <= IO_9_5_IN_pin_0_driver_mux_fanins(IO_9_5_IN_pin_0_driver_mux_selector);
	IO_9_5_IN_pin_1  <= IO_9_5_IN_pin_1_driver_mux_fanins(IO_9_5_IN_pin_1_driver_mux_selector);
	IO_9_6_IN_pin_0  <= IO_9_6_IN_pin_0_driver_mux_fanins(IO_9_6_IN_pin_0_driver_mux_selector);
	IO_9_6_IN_pin_1  <= IO_9_6_IN_pin_1_driver_mux_fanins(IO_9_6_IN_pin_1_driver_mux_selector);

	-- Tracks fanin choices (inputs of the mux driving the track) --
	track_0_1_chanY_n0_driver_mux_fanins  <= "0" & IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_0_chanX_n3;
	track_0_1_chanY_n1_driver_mux_fanins  <= IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_1_chanX_n1 & track_0_2_chanY_n1;
	track_0_1_chanY_n10_driver_mux_fanins <= IO_0_1_OUT_pin_1 & track_1_0_chanX_n13;
	track_0_1_chanY_n11_driver_mux_fanins <= "0" & IO_0_1_OUT_pin_1 & track_1_1_chanX_n11 & track_0_2_chanY_n11;
	track_0_1_chanY_n12_driver_mux_fanins <= IO_0_1_OUT_pin_1 & track_1_0_chanX_n15;
	track_0_1_chanY_n13_driver_mux_fanins <= "0" & IO_0_1_OUT_pin_1 & track_1_1_chanX_n13 & track_0_2_chanY_n13;
	track_0_1_chanY_n14_driver_mux_fanins <= IO_0_1_OUT_pin_1 & track_1_0_chanX_n1;
	track_0_1_chanY_n15_driver_mux_fanins <= "0" & IO_0_1_OUT_pin_1 & track_1_1_chanX_n15 & track_0_2_chanY_n15;
	track_0_1_chanY_n2_driver_mux_fanins  <= "0" & IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_0_chanX_n5;
	track_0_1_chanY_n3_driver_mux_fanins  <= IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_1_chanX_n3 & track_0_2_chanY_n3;
	track_0_1_chanY_n4_driver_mux_fanins  <= "0" & IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_0_chanX_n7;
	track_0_1_chanY_n5_driver_mux_fanins  <= IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_1_chanX_n5 & track_0_2_chanY_n5;
	track_0_1_chanY_n6_driver_mux_fanins  <= "0" & IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_0_chanX_n9;
	track_0_1_chanY_n7_driver_mux_fanins  <= IO_0_1_OUT_pin_0 & CLB_1_1_OUT_pin_1 & track_1_1_chanX_n7 & track_0_2_chanY_n7;
	track_0_1_chanY_n8_driver_mux_fanins  <= IO_0_1_OUT_pin_1 & track_1_0_chanX_n11;
	track_0_1_chanY_n9_driver_mux_fanins  <= "0" & IO_0_1_OUT_pin_1 & track_1_1_chanX_n9 & track_0_2_chanY_n9;
	track_0_2_chanY_n0_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_0_1_chanY_n0 & track_1_1_chanX_n1;
	track_0_2_chanY_n1_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_1_2_chanX_n1 & track_0_3_chanY_n1;
	track_0_2_chanY_n10_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_0_1_chanY_n10 & track_1_1_chanX_n11;
	track_0_2_chanY_n11_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_1_2_chanX_n11 & track_0_3_chanY_n11;
	track_0_2_chanY_n12_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_0_1_chanY_n12 & track_1_1_chanX_n13;
	track_0_2_chanY_n13_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_1_2_chanX_n13 & track_0_3_chanY_n13;
	track_0_2_chanY_n14_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_0_1_chanY_n14 & track_1_1_chanX_n15;
	track_0_2_chanY_n15_driver_mux_fanins <= "0" & IO_0_2_OUT_pin_1 & track_1_2_chanX_n15 & track_0_3_chanY_n15;
	track_0_2_chanY_n2_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_0_1_chanY_n2 & track_1_1_chanX_n3;
	track_0_2_chanY_n3_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_1_2_chanX_n3 & track_0_3_chanY_n3;
	track_0_2_chanY_n4_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_0_1_chanY_n4 & track_1_1_chanX_n5;
	track_0_2_chanY_n5_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_1_2_chanX_n5 & track_0_3_chanY_n5;
	track_0_2_chanY_n6_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_0_1_chanY_n6 & track_1_1_chanX_n7;
	track_0_2_chanY_n7_driver_mux_fanins  <= IO_0_2_OUT_pin_0 & CLB_1_2_OUT_pin_1 & track_1_2_chanX_n7 & track_0_3_chanY_n7;
	track_0_2_chanY_n8_driver_mux_fanins  <= "0" & IO_0_2_OUT_pin_1 & track_0_1_chanY_n8 & track_1_1_chanX_n9;
	track_0_2_chanY_n9_driver_mux_fanins  <= "0" & IO_0_2_OUT_pin_1 & track_1_2_chanX_n9 & track_0_3_chanY_n9;
	track_0_3_chanY_n0_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_0_2_chanY_n0 & track_1_2_chanX_n1;
	track_0_3_chanY_n1_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_1_3_chanX_n1 & track_0_4_chanY_n1;
	track_0_3_chanY_n10_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_0_2_chanY_n10 & track_1_2_chanX_n11;
	track_0_3_chanY_n11_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_1_3_chanX_n11 & track_0_4_chanY_n11;
	track_0_3_chanY_n12_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_0_2_chanY_n12 & track_1_2_chanX_n13;
	track_0_3_chanY_n13_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_1_3_chanX_n13 & track_0_4_chanY_n13;
	track_0_3_chanY_n14_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_0_2_chanY_n14 & track_1_2_chanX_n15;
	track_0_3_chanY_n15_driver_mux_fanins <= "0" & IO_0_3_OUT_pin_1 & track_1_3_chanX_n15 & track_0_4_chanY_n15;
	track_0_3_chanY_n2_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_0_2_chanY_n2 & track_1_2_chanX_n3;
	track_0_3_chanY_n3_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_1_3_chanX_n3 & track_0_4_chanY_n3;
	track_0_3_chanY_n4_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_0_2_chanY_n4 & track_1_2_chanX_n5;
	track_0_3_chanY_n5_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_1_3_chanX_n5 & track_0_4_chanY_n5;
	track_0_3_chanY_n6_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_0_2_chanY_n6 & track_1_2_chanX_n7;
	track_0_3_chanY_n7_driver_mux_fanins  <= IO_0_3_OUT_pin_0 & CLB_1_3_OUT_pin_1 & track_1_3_chanX_n7 & track_0_4_chanY_n7;
	track_0_3_chanY_n8_driver_mux_fanins  <= "0" & IO_0_3_OUT_pin_1 & track_0_2_chanY_n8 & track_1_2_chanX_n9;
	track_0_3_chanY_n9_driver_mux_fanins  <= "0" & IO_0_3_OUT_pin_1 & track_1_3_chanX_n9 & track_0_4_chanY_n9;
	track_0_4_chanY_n0_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_0_3_chanY_n0 & track_1_3_chanX_n1;
	track_0_4_chanY_n1_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_1_4_chanX_n1 & track_0_5_chanY_n1;
	track_0_4_chanY_n10_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_0_3_chanY_n10 & track_1_3_chanX_n11;
	track_0_4_chanY_n11_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_1_4_chanX_n11 & track_0_5_chanY_n11;
	track_0_4_chanY_n12_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_0_3_chanY_n12 & track_1_3_chanX_n13;
	track_0_4_chanY_n13_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_1_4_chanX_n13 & track_0_5_chanY_n13;
	track_0_4_chanY_n14_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_0_3_chanY_n14 & track_1_3_chanX_n15;
	track_0_4_chanY_n15_driver_mux_fanins <= "0" & IO_0_4_OUT_pin_1 & track_1_4_chanX_n15 & track_0_5_chanY_n15;
	track_0_4_chanY_n2_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_0_3_chanY_n2 & track_1_3_chanX_n3;
	track_0_4_chanY_n3_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_1_4_chanX_n3 & track_0_5_chanY_n3;
	track_0_4_chanY_n4_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_0_3_chanY_n4 & track_1_3_chanX_n5;
	track_0_4_chanY_n5_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_1_4_chanX_n5 & track_0_5_chanY_n5;
	track_0_4_chanY_n6_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_0_3_chanY_n6 & track_1_3_chanX_n7;
	track_0_4_chanY_n7_driver_mux_fanins  <= IO_0_4_OUT_pin_0 & CLB_1_4_OUT_pin_1 & track_1_4_chanX_n7 & track_0_5_chanY_n7;
	track_0_4_chanY_n8_driver_mux_fanins  <= "0" & IO_0_4_OUT_pin_1 & track_0_3_chanY_n8 & track_1_3_chanX_n9;
	track_0_4_chanY_n9_driver_mux_fanins  <= "0" & IO_0_4_OUT_pin_1 & track_1_4_chanX_n9 & track_0_5_chanY_n9;
	track_0_5_chanY_n0_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_0_4_chanY_n0 & track_1_4_chanX_n1;
	track_0_5_chanY_n1_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_1_5_chanX_n1 & track_0_6_chanY_n1;
	track_0_5_chanY_n10_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_0_4_chanY_n10 & track_1_4_chanX_n11;
	track_0_5_chanY_n11_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_1_5_chanX_n11 & track_0_6_chanY_n11;
	track_0_5_chanY_n12_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_0_4_chanY_n12 & track_1_4_chanX_n13;
	track_0_5_chanY_n13_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_1_5_chanX_n13 & track_0_6_chanY_n13;
	track_0_5_chanY_n14_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_0_4_chanY_n14 & track_1_4_chanX_n15;
	track_0_5_chanY_n15_driver_mux_fanins <= "0" & IO_0_5_OUT_pin_1 & track_1_5_chanX_n15 & track_0_6_chanY_n15;
	track_0_5_chanY_n2_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_0_4_chanY_n2 & track_1_4_chanX_n3;
	track_0_5_chanY_n3_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_1_5_chanX_n3 & track_0_6_chanY_n3;
	track_0_5_chanY_n4_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_0_4_chanY_n4 & track_1_4_chanX_n5;
	track_0_5_chanY_n5_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_1_5_chanX_n5 & track_0_6_chanY_n5;
	track_0_5_chanY_n6_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_0_4_chanY_n6 & track_1_4_chanX_n7;
	track_0_5_chanY_n7_driver_mux_fanins  <= IO_0_5_OUT_pin_0 & CLB_1_5_OUT_pin_1 & track_1_5_chanX_n7 & track_0_6_chanY_n7;
	track_0_5_chanY_n8_driver_mux_fanins  <= "0" & IO_0_5_OUT_pin_1 & track_0_4_chanY_n8 & track_1_4_chanX_n9;
	track_0_5_chanY_n9_driver_mux_fanins  <= "0" & IO_0_5_OUT_pin_1 & track_1_5_chanX_n9 & track_0_6_chanY_n9;
	track_0_6_chanY_n0_driver_mux_fanins  <= IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_0_5_chanY_n0 & track_1_5_chanX_n1;
	track_0_6_chanY_n1_driver_mux_fanins  <= "0" & IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_1_6_chanX_n13;
	track_0_6_chanY_n10_driver_mux_fanins <= "0" & IO_0_6_OUT_pin_1 & track_0_5_chanY_n10 & track_1_5_chanX_n11;
	track_0_6_chanY_n11_driver_mux_fanins <= IO_0_6_OUT_pin_1 & track_1_6_chanX_n3;
	track_0_6_chanY_n12_driver_mux_fanins <= "0" & IO_0_6_OUT_pin_1 & track_0_5_chanY_n12 & track_1_5_chanX_n13;
	track_0_6_chanY_n13_driver_mux_fanins <= IO_0_6_OUT_pin_1 & track_1_6_chanX_n1;
	track_0_6_chanY_n14_driver_mux_fanins <= "0" & IO_0_6_OUT_pin_1 & track_0_5_chanY_n14 & track_1_5_chanX_n15;
	track_0_6_chanY_n15_driver_mux_fanins <= IO_0_6_OUT_pin_1 & track_1_6_chanX_n15;
	track_0_6_chanY_n2_driver_mux_fanins  <= IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_0_5_chanY_n2 & track_1_5_chanX_n3;
	track_0_6_chanY_n3_driver_mux_fanins  <= "0" & IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_1_6_chanX_n11;
	track_0_6_chanY_n4_driver_mux_fanins  <= IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_0_5_chanY_n4 & track_1_5_chanX_n5;
	track_0_6_chanY_n5_driver_mux_fanins  <= "0" & IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_1_6_chanX_n9;
	track_0_6_chanY_n6_driver_mux_fanins  <= IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_0_5_chanY_n6 & track_1_5_chanX_n7;
	track_0_6_chanY_n7_driver_mux_fanins  <= "0" & IO_0_6_OUT_pin_0 & CLB_1_6_OUT_pin_1 & track_1_6_chanX_n7;
	track_0_6_chanY_n8_driver_mux_fanins  <= "0" & IO_0_6_OUT_pin_1 & track_0_5_chanY_n8 & track_1_5_chanX_n9;
	track_0_6_chanY_n9_driver_mux_fanins  <= IO_0_6_OUT_pin_1 & track_1_6_chanX_n5;
	track_1_0_chanX_n0_driver_mux_fanins  <= "0" & IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_0_1_chanY_n15;
	track_1_0_chanX_n1_driver_mux_fanins  <= IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_2_0_chanX_n1 & track_1_1_chanY_n1;
	track_1_0_chanX_n10_driver_mux_fanins <= IO_1_0_OUT_pin_1 & track_0_1_chanY_n9;
	track_1_0_chanX_n11_driver_mux_fanins <= "0" & IO_1_0_OUT_pin_1 & track_2_0_chanX_n11 & track_1_1_chanY_n11;
	track_1_0_chanX_n12_driver_mux_fanins <= IO_1_0_OUT_pin_1 & track_0_1_chanY_n11;
	track_1_0_chanX_n13_driver_mux_fanins <= "0" & IO_1_0_OUT_pin_1 & track_2_0_chanX_n13 & track_1_1_chanY_n13;
	track_1_0_chanX_n14_driver_mux_fanins <= IO_1_0_OUT_pin_1 & track_0_1_chanY_n13;
	track_1_0_chanX_n15_driver_mux_fanins <= "0" & IO_1_0_OUT_pin_1 & track_2_0_chanX_n15 & track_1_1_chanY_n15;
	track_1_0_chanX_n2_driver_mux_fanins  <= "0" & IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_0_1_chanY_n1;
	track_1_0_chanX_n3_driver_mux_fanins  <= IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_2_0_chanX_n3 & track_1_1_chanY_n3;
	track_1_0_chanX_n4_driver_mux_fanins  <= "0" & IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_0_1_chanY_n3;
	track_1_0_chanX_n5_driver_mux_fanins  <= IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_2_0_chanX_n5 & track_1_1_chanY_n5;
	track_1_0_chanX_n6_driver_mux_fanins  <= "0" & IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_0_1_chanY_n5;
	track_1_0_chanX_n7_driver_mux_fanins  <= IO_1_0_OUT_pin_0 & CLB_1_1_OUT_pin_0 & track_2_0_chanX_n7 & track_1_1_chanY_n7;
	track_1_0_chanX_n8_driver_mux_fanins  <= IO_1_0_OUT_pin_1 & track_0_1_chanY_n7;
	track_1_0_chanX_n9_driver_mux_fanins  <= "0" & IO_1_0_OUT_pin_1 & track_2_0_chanX_n9 & track_1_1_chanY_n9;
	track_1_1_chanX_n0_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_2 & track_0_1_chanY_n6 & track_0_2_chanY_n7;
	track_1_1_chanX_n1_driver_mux_fanins  <= CLB_1_1_OUT_pin_2 & track_1_1_chanY_n14 & track_2_1_chanX_n1 & track_1_2_chanY_n1;
	track_1_1_chanX_n10_driver_mux_fanins <= "0" & CLB_1_2_OUT_pin_0 & track_0_1_chanY_n10 & track_0_2_chanY_n11;
	track_1_1_chanX_n11_driver_mux_fanins <= CLB_1_2_OUT_pin_0 & track_1_1_chanY_n8 & track_2_1_chanX_n11 & track_1_2_chanY_n7;
	track_1_1_chanX_n12_driver_mux_fanins <= "0" & CLB_1_2_OUT_pin_0 & track_0_1_chanY_n12 & track_0_2_chanY_n13;
	track_1_1_chanX_n13_driver_mux_fanins <= CLB_1_2_OUT_pin_0 & track_1_1_chanY_n10 & track_2_1_chanX_n13 & track_1_2_chanY_n5;
	track_1_1_chanX_n14_driver_mux_fanins <= "0" & CLB_1_2_OUT_pin_0 & track_0_1_chanY_n14 & track_0_2_chanY_n15;
	track_1_1_chanX_n15_driver_mux_fanins <= CLB_1_2_OUT_pin_0 & track_1_1_chanY_n12 & track_2_1_chanX_n15 & track_1_2_chanY_n3;
	track_1_1_chanX_n2_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_2 & track_0_1_chanY_n8 & track_0_2_chanY_n9;
	track_1_1_chanX_n3_driver_mux_fanins  <= CLB_1_1_OUT_pin_2 & track_1_1_chanY_n0 & track_2_1_chanX_n3 & track_1_2_chanY_n15;
	track_1_1_chanX_n4_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_2 & track_0_1_chanY_n0 & track_0_2_chanY_n1;
	track_1_1_chanX_n5_driver_mux_fanins  <= CLB_1_1_OUT_pin_2 & track_1_1_chanY_n2 & track_2_1_chanX_n5 & track_1_2_chanY_n13;
	track_1_1_chanX_n6_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_2 & track_0_1_chanY_n2 & track_0_2_chanY_n3;
	track_1_1_chanX_n7_driver_mux_fanins  <= CLB_1_1_OUT_pin_2 & track_1_1_chanY_n4 & track_2_1_chanX_n7 & track_1_2_chanY_n11;
	track_1_1_chanX_n8_driver_mux_fanins  <= "0" & CLB_1_2_OUT_pin_0 & track_0_1_chanY_n4 & track_0_2_chanY_n5;
	track_1_1_chanX_n9_driver_mux_fanins  <= CLB_1_2_OUT_pin_0 & track_1_1_chanY_n6 & track_2_1_chanX_n9 & track_1_2_chanY_n9;
	track_1_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_3 & track_2_0_chanX_n7 & track_1_0_chanX_n6;
	track_1_1_chanY_n1_driver_mux_fanins  <= CLB_1_1_OUT_pin_3 & track_2_1_chanX_n13 & track_1_1_chanX_n2 & track_1_2_chanY_n1;
	track_1_1_chanY_n10_driver_mux_fanins <= "0" & CLB_2_1_OUT_pin_1 & track_2_0_chanX_n11 & track_1_0_chanX_n10;
	track_1_1_chanY_n11_driver_mux_fanins <= CLB_2_1_OUT_pin_1 & track_2_1_chanX_n3 & track_1_1_chanX_n12 & track_1_2_chanY_n11;
	track_1_1_chanY_n12_driver_mux_fanins <= "0" & CLB_2_1_OUT_pin_1 & track_2_0_chanX_n13 & track_1_0_chanX_n12;
	track_1_1_chanY_n13_driver_mux_fanins <= CLB_2_1_OUT_pin_1 & track_2_1_chanX_n1 & track_1_1_chanX_n14 & track_1_2_chanY_n13;
	track_1_1_chanY_n14_driver_mux_fanins <= "0" & CLB_2_1_OUT_pin_1 & track_2_0_chanX_n15 & track_1_0_chanX_n14;
	track_1_1_chanY_n15_driver_mux_fanins <= CLB_2_1_OUT_pin_1 & track_2_1_chanX_n15 & track_1_1_chanX_n0 & track_1_2_chanY_n15;
	track_1_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_3 & track_2_0_chanX_n9 & track_1_0_chanX_n8;
	track_1_1_chanY_n3_driver_mux_fanins  <= CLB_1_1_OUT_pin_3 & track_2_1_chanX_n11 & track_1_1_chanX_n4 & track_1_2_chanY_n3;
	track_1_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_3 & track_2_0_chanX_n1 & track_1_0_chanX_n0;
	track_1_1_chanY_n5_driver_mux_fanins  <= CLB_1_1_OUT_pin_3 & track_2_1_chanX_n9 & track_1_1_chanX_n6 & track_1_2_chanY_n5;
	track_1_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_1_1_OUT_pin_3 & track_2_0_chanX_n3 & track_1_0_chanX_n2;
	track_1_1_chanY_n7_driver_mux_fanins  <= CLB_1_1_OUT_pin_3 & track_2_1_chanX_n7 & track_1_1_chanX_n8 & track_1_2_chanY_n7;
	track_1_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_2_1_OUT_pin_1 & track_2_0_chanX_n5 & track_1_0_chanX_n4;
	track_1_1_chanY_n9_driver_mux_fanins  <= CLB_2_1_OUT_pin_1 & track_2_1_chanX_n5 & track_1_1_chanX_n10 & track_1_2_chanY_n9;
	track_1_2_chanX_n0_driver_mux_fanins  <= "0" & CLB_1_2_OUT_pin_2 & track_0_2_chanY_n6 & track_0_3_chanY_n7;
	track_1_2_chanX_n1_driver_mux_fanins  <= CLB_1_2_OUT_pin_2 & track_1_2_chanY_n14 & track_2_2_chanX_n1 & track_1_3_chanY_n1;
	track_1_2_chanX_n10_driver_mux_fanins <= "0" & CLB_1_3_OUT_pin_0 & track_0_2_chanY_n10 & track_0_3_chanY_n11;
	track_1_2_chanX_n11_driver_mux_fanins <= CLB_1_3_OUT_pin_0 & track_1_2_chanY_n8 & track_2_2_chanX_n11 & track_1_3_chanY_n7;
	track_1_2_chanX_n12_driver_mux_fanins <= "0" & CLB_1_3_OUT_pin_0 & track_0_2_chanY_n12 & track_0_3_chanY_n13;
	track_1_2_chanX_n13_driver_mux_fanins <= CLB_1_3_OUT_pin_0 & track_1_2_chanY_n10 & track_2_2_chanX_n13 & track_1_3_chanY_n5;
	track_1_2_chanX_n14_driver_mux_fanins <= "0" & CLB_1_3_OUT_pin_0 & track_0_2_chanY_n14 & track_0_3_chanY_n15;
	track_1_2_chanX_n15_driver_mux_fanins <= CLB_1_3_OUT_pin_0 & track_1_2_chanY_n12 & track_2_2_chanX_n15 & track_1_3_chanY_n3;
	track_1_2_chanX_n2_driver_mux_fanins  <= "0" & CLB_1_2_OUT_pin_2 & track_0_2_chanY_n8 & track_0_3_chanY_n9;
	track_1_2_chanX_n3_driver_mux_fanins  <= CLB_1_2_OUT_pin_2 & track_1_2_chanY_n0 & track_2_2_chanX_n3 & track_1_3_chanY_n15;
	track_1_2_chanX_n4_driver_mux_fanins  <= "0" & CLB_1_2_OUT_pin_2 & track_0_2_chanY_n0 & track_0_3_chanY_n1;
	track_1_2_chanX_n5_driver_mux_fanins  <= CLB_1_2_OUT_pin_2 & track_1_2_chanY_n2 & track_2_2_chanX_n5 & track_1_3_chanY_n13;
	track_1_2_chanX_n6_driver_mux_fanins  <= "0" & CLB_1_2_OUT_pin_2 & track_0_2_chanY_n2 & track_0_3_chanY_n3;
	track_1_2_chanX_n7_driver_mux_fanins  <= CLB_1_2_OUT_pin_2 & track_1_2_chanY_n4 & track_2_2_chanX_n7 & track_1_3_chanY_n11;
	track_1_2_chanX_n8_driver_mux_fanins  <= "0" & CLB_1_3_OUT_pin_0 & track_0_2_chanY_n4 & track_0_3_chanY_n5;
	track_1_2_chanX_n9_driver_mux_fanins  <= CLB_1_3_OUT_pin_0 & track_1_2_chanY_n6 & track_2_2_chanX_n9 & track_1_3_chanY_n9;
	track_1_2_chanY_n0_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_1_1_chanY_n0 & track_2_1_chanX_n3 & track_1_1_chanX_n0;
	track_1_2_chanY_n1_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_2_2_chanX_n13 & track_1_2_chanX_n2 & track_1_3_chanY_n1;
	track_1_2_chanY_n10_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_1_1_chanY_n10 & track_2_1_chanX_n13 & track_1_1_chanX_n6;
	track_1_2_chanY_n11_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_2_2_chanX_n3 & track_1_2_chanX_n12 & track_1_3_chanY_n11;
	track_1_2_chanY_n12_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_1_1_chanY_n12 & track_2_1_chanX_n15 & track_1_1_chanX_n4;
	track_1_2_chanY_n13_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_2_2_chanX_n1 & track_1_2_chanX_n14 & track_1_3_chanY_n13;
	track_1_2_chanY_n14_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_1_1_chanY_n14 & track_2_1_chanX_n1 & track_1_1_chanX_n2;
	track_1_2_chanY_n15_driver_mux_fanins <= CLB_2_2_OUT_pin_1 & track_2_2_chanX_n15 & track_1_2_chanX_n0 & track_1_3_chanY_n15;
	track_1_2_chanY_n2_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_1_1_chanY_n2 & track_2_1_chanX_n5 & track_1_1_chanX_n14;
	track_1_2_chanY_n3_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_2_2_chanX_n11 & track_1_2_chanX_n4 & track_1_3_chanY_n3;
	track_1_2_chanY_n4_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_1_1_chanY_n4 & track_2_1_chanX_n7 & track_1_1_chanX_n12;
	track_1_2_chanY_n5_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_2_2_chanX_n9 & track_1_2_chanX_n6 & track_1_3_chanY_n5;
	track_1_2_chanY_n6_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_1_1_chanY_n6 & track_2_1_chanX_n9 & track_1_1_chanX_n10;
	track_1_2_chanY_n7_driver_mux_fanins  <= CLB_1_2_OUT_pin_3 & track_2_2_chanX_n7 & track_1_2_chanX_n8 & track_1_3_chanY_n7;
	track_1_2_chanY_n8_driver_mux_fanins  <= CLB_2_2_OUT_pin_1 & track_1_1_chanY_n8 & track_2_1_chanX_n11 & track_1_1_chanX_n8;
	track_1_2_chanY_n9_driver_mux_fanins  <= CLB_2_2_OUT_pin_1 & track_2_2_chanX_n5 & track_1_2_chanX_n10 & track_1_3_chanY_n9;
	track_1_3_chanX_n0_driver_mux_fanins  <= "0" & CLB_1_3_OUT_pin_2 & track_0_3_chanY_n6 & track_0_4_chanY_n7;
	track_1_3_chanX_n1_driver_mux_fanins  <= CLB_1_3_OUT_pin_2 & track_1_3_chanY_n14 & track_2_3_chanX_n1 & track_1_4_chanY_n1;
	track_1_3_chanX_n10_driver_mux_fanins <= "0" & CLB_1_4_OUT_pin_0 & track_0_3_chanY_n10 & track_0_4_chanY_n11;
	track_1_3_chanX_n11_driver_mux_fanins <= CLB_1_4_OUT_pin_0 & track_1_3_chanY_n8 & track_2_3_chanX_n11 & track_1_4_chanY_n7;
	track_1_3_chanX_n12_driver_mux_fanins <= "0" & CLB_1_4_OUT_pin_0 & track_0_3_chanY_n12 & track_0_4_chanY_n13;
	track_1_3_chanX_n13_driver_mux_fanins <= CLB_1_4_OUT_pin_0 & track_1_3_chanY_n10 & track_2_3_chanX_n13 & track_1_4_chanY_n5;
	track_1_3_chanX_n14_driver_mux_fanins <= "0" & CLB_1_4_OUT_pin_0 & track_0_3_chanY_n14 & track_0_4_chanY_n15;
	track_1_3_chanX_n15_driver_mux_fanins <= CLB_1_4_OUT_pin_0 & track_1_3_chanY_n12 & track_2_3_chanX_n15 & track_1_4_chanY_n3;
	track_1_3_chanX_n2_driver_mux_fanins  <= "0" & CLB_1_3_OUT_pin_2 & track_0_3_chanY_n8 & track_0_4_chanY_n9;
	track_1_3_chanX_n3_driver_mux_fanins  <= CLB_1_3_OUT_pin_2 & track_1_3_chanY_n0 & track_2_3_chanX_n3 & track_1_4_chanY_n15;
	track_1_3_chanX_n4_driver_mux_fanins  <= "0" & CLB_1_3_OUT_pin_2 & track_0_3_chanY_n0 & track_0_4_chanY_n1;
	track_1_3_chanX_n5_driver_mux_fanins  <= CLB_1_3_OUT_pin_2 & track_1_3_chanY_n2 & track_2_3_chanX_n5 & track_1_4_chanY_n13;
	track_1_3_chanX_n6_driver_mux_fanins  <= "0" & CLB_1_3_OUT_pin_2 & track_0_3_chanY_n2 & track_0_4_chanY_n3;
	track_1_3_chanX_n7_driver_mux_fanins  <= CLB_1_3_OUT_pin_2 & track_1_3_chanY_n4 & track_2_3_chanX_n7 & track_1_4_chanY_n11;
	track_1_3_chanX_n8_driver_mux_fanins  <= "0" & CLB_1_4_OUT_pin_0 & track_0_3_chanY_n4 & track_0_4_chanY_n5;
	track_1_3_chanX_n9_driver_mux_fanins  <= CLB_1_4_OUT_pin_0 & track_1_3_chanY_n6 & track_2_3_chanX_n9 & track_1_4_chanY_n9;
	track_1_3_chanY_n0_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_1_2_chanY_n0 & track_2_2_chanX_n3 & track_1_2_chanX_n0;
	track_1_3_chanY_n1_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_2_3_chanX_n13 & track_1_3_chanX_n2 & track_1_4_chanY_n1;
	track_1_3_chanY_n10_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_1_2_chanY_n10 & track_2_2_chanX_n13 & track_1_2_chanX_n6;
	track_1_3_chanY_n11_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_2_3_chanX_n3 & track_1_3_chanX_n12 & track_1_4_chanY_n11;
	track_1_3_chanY_n12_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_1_2_chanY_n12 & track_2_2_chanX_n15 & track_1_2_chanX_n4;
	track_1_3_chanY_n13_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_2_3_chanX_n1 & track_1_3_chanX_n14 & track_1_4_chanY_n13;
	track_1_3_chanY_n14_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_1_2_chanY_n14 & track_2_2_chanX_n1 & track_1_2_chanX_n2;
	track_1_3_chanY_n15_driver_mux_fanins <= CLB_2_3_OUT_pin_1 & track_2_3_chanX_n15 & track_1_3_chanX_n0 & track_1_4_chanY_n15;
	track_1_3_chanY_n2_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_1_2_chanY_n2 & track_2_2_chanX_n5 & track_1_2_chanX_n14;
	track_1_3_chanY_n3_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_2_3_chanX_n11 & track_1_3_chanX_n4 & track_1_4_chanY_n3;
	track_1_3_chanY_n4_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_1_2_chanY_n4 & track_2_2_chanX_n7 & track_1_2_chanX_n12;
	track_1_3_chanY_n5_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_2_3_chanX_n9 & track_1_3_chanX_n6 & track_1_4_chanY_n5;
	track_1_3_chanY_n6_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_1_2_chanY_n6 & track_2_2_chanX_n9 & track_1_2_chanX_n10;
	track_1_3_chanY_n7_driver_mux_fanins  <= CLB_1_3_OUT_pin_3 & track_2_3_chanX_n7 & track_1_3_chanX_n8 & track_1_4_chanY_n7;
	track_1_3_chanY_n8_driver_mux_fanins  <= CLB_2_3_OUT_pin_1 & track_1_2_chanY_n8 & track_2_2_chanX_n11 & track_1_2_chanX_n8;
	track_1_3_chanY_n9_driver_mux_fanins  <= CLB_2_3_OUT_pin_1 & track_2_3_chanX_n5 & track_1_3_chanX_n10 & track_1_4_chanY_n9;
	track_1_4_chanX_n0_driver_mux_fanins  <= "0" & CLB_1_4_OUT_pin_2 & track_0_4_chanY_n6 & track_0_5_chanY_n7;
	track_1_4_chanX_n1_driver_mux_fanins  <= CLB_1_4_OUT_pin_2 & track_1_4_chanY_n14 & track_2_4_chanX_n1 & track_1_5_chanY_n1;
	track_1_4_chanX_n10_driver_mux_fanins <= "0" & CLB_1_5_OUT_pin_0 & track_0_4_chanY_n10 & track_0_5_chanY_n11;
	track_1_4_chanX_n11_driver_mux_fanins <= CLB_1_5_OUT_pin_0 & track_1_4_chanY_n8 & track_2_4_chanX_n11 & track_1_5_chanY_n7;
	track_1_4_chanX_n12_driver_mux_fanins <= "0" & CLB_1_5_OUT_pin_0 & track_0_4_chanY_n12 & track_0_5_chanY_n13;
	track_1_4_chanX_n13_driver_mux_fanins <= CLB_1_5_OUT_pin_0 & track_1_4_chanY_n10 & track_2_4_chanX_n13 & track_1_5_chanY_n5;
	track_1_4_chanX_n14_driver_mux_fanins <= "0" & CLB_1_5_OUT_pin_0 & track_0_4_chanY_n14 & track_0_5_chanY_n15;
	track_1_4_chanX_n15_driver_mux_fanins <= CLB_1_5_OUT_pin_0 & track_1_4_chanY_n12 & track_2_4_chanX_n15 & track_1_5_chanY_n3;
	track_1_4_chanX_n2_driver_mux_fanins  <= "0" & CLB_1_4_OUT_pin_2 & track_0_4_chanY_n8 & track_0_5_chanY_n9;
	track_1_4_chanX_n3_driver_mux_fanins  <= CLB_1_4_OUT_pin_2 & track_1_4_chanY_n0 & track_2_4_chanX_n3 & track_1_5_chanY_n15;
	track_1_4_chanX_n4_driver_mux_fanins  <= "0" & CLB_1_4_OUT_pin_2 & track_0_4_chanY_n0 & track_0_5_chanY_n1;
	track_1_4_chanX_n5_driver_mux_fanins  <= CLB_1_4_OUT_pin_2 & track_1_4_chanY_n2 & track_2_4_chanX_n5 & track_1_5_chanY_n13;
	track_1_4_chanX_n6_driver_mux_fanins  <= "0" & CLB_1_4_OUT_pin_2 & track_0_4_chanY_n2 & track_0_5_chanY_n3;
	track_1_4_chanX_n7_driver_mux_fanins  <= CLB_1_4_OUT_pin_2 & track_1_4_chanY_n4 & track_2_4_chanX_n7 & track_1_5_chanY_n11;
	track_1_4_chanX_n8_driver_mux_fanins  <= "0" & CLB_1_5_OUT_pin_0 & track_0_4_chanY_n4 & track_0_5_chanY_n5;
	track_1_4_chanX_n9_driver_mux_fanins  <= CLB_1_5_OUT_pin_0 & track_1_4_chanY_n6 & track_2_4_chanX_n9 & track_1_5_chanY_n9;
	track_1_4_chanY_n0_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_1_3_chanY_n0 & track_2_3_chanX_n3 & track_1_3_chanX_n0;
	track_1_4_chanY_n1_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_2_4_chanX_n13 & track_1_4_chanX_n2 & track_1_5_chanY_n1;
	track_1_4_chanY_n10_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_1_3_chanY_n10 & track_2_3_chanX_n13 & track_1_3_chanX_n6;
	track_1_4_chanY_n11_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_2_4_chanX_n3 & track_1_4_chanX_n12 & track_1_5_chanY_n11;
	track_1_4_chanY_n12_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_1_3_chanY_n12 & track_2_3_chanX_n15 & track_1_3_chanX_n4;
	track_1_4_chanY_n13_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_2_4_chanX_n1 & track_1_4_chanX_n14 & track_1_5_chanY_n13;
	track_1_4_chanY_n14_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_1_3_chanY_n14 & track_2_3_chanX_n1 & track_1_3_chanX_n2;
	track_1_4_chanY_n15_driver_mux_fanins <= CLB_2_4_OUT_pin_1 & track_2_4_chanX_n15 & track_1_4_chanX_n0 & track_1_5_chanY_n15;
	track_1_4_chanY_n2_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_1_3_chanY_n2 & track_2_3_chanX_n5 & track_1_3_chanX_n14;
	track_1_4_chanY_n3_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_2_4_chanX_n11 & track_1_4_chanX_n4 & track_1_5_chanY_n3;
	track_1_4_chanY_n4_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_1_3_chanY_n4 & track_2_3_chanX_n7 & track_1_3_chanX_n12;
	track_1_4_chanY_n5_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_2_4_chanX_n9 & track_1_4_chanX_n6 & track_1_5_chanY_n5;
	track_1_4_chanY_n6_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_1_3_chanY_n6 & track_2_3_chanX_n9 & track_1_3_chanX_n10;
	track_1_4_chanY_n7_driver_mux_fanins  <= CLB_1_4_OUT_pin_3 & track_2_4_chanX_n7 & track_1_4_chanX_n8 & track_1_5_chanY_n7;
	track_1_4_chanY_n8_driver_mux_fanins  <= CLB_2_4_OUT_pin_1 & track_1_3_chanY_n8 & track_2_3_chanX_n11 & track_1_3_chanX_n8;
	track_1_4_chanY_n9_driver_mux_fanins  <= CLB_2_4_OUT_pin_1 & track_2_4_chanX_n5 & track_1_4_chanX_n10 & track_1_5_chanY_n9;
	track_1_5_chanX_n0_driver_mux_fanins  <= "0" & CLB_1_5_OUT_pin_2 & track_0_5_chanY_n6 & track_0_6_chanY_n7;
	track_1_5_chanX_n1_driver_mux_fanins  <= CLB_1_5_OUT_pin_2 & track_1_5_chanY_n14 & track_2_5_chanX_n1 & track_1_6_chanY_n1;
	track_1_5_chanX_n10_driver_mux_fanins <= "0" & CLB_1_6_OUT_pin_0 & track_0_5_chanY_n10 & track_0_6_chanY_n11;
	track_1_5_chanX_n11_driver_mux_fanins <= CLB_1_6_OUT_pin_0 & track_1_5_chanY_n8 & track_2_5_chanX_n11 & track_1_6_chanY_n7;
	track_1_5_chanX_n12_driver_mux_fanins <= "0" & CLB_1_6_OUT_pin_0 & track_0_5_chanY_n12 & track_0_6_chanY_n13;
	track_1_5_chanX_n13_driver_mux_fanins <= CLB_1_6_OUT_pin_0 & track_1_5_chanY_n10 & track_2_5_chanX_n13 & track_1_6_chanY_n5;
	track_1_5_chanX_n14_driver_mux_fanins <= "0" & CLB_1_6_OUT_pin_0 & track_0_5_chanY_n14 & track_0_6_chanY_n15;
	track_1_5_chanX_n15_driver_mux_fanins <= CLB_1_6_OUT_pin_0 & track_1_5_chanY_n12 & track_2_5_chanX_n15 & track_1_6_chanY_n3;
	track_1_5_chanX_n2_driver_mux_fanins  <= "0" & CLB_1_5_OUT_pin_2 & track_0_5_chanY_n8 & track_0_6_chanY_n9;
	track_1_5_chanX_n3_driver_mux_fanins  <= CLB_1_5_OUT_pin_2 & track_1_5_chanY_n0 & track_2_5_chanX_n3 & track_1_6_chanY_n15;
	track_1_5_chanX_n4_driver_mux_fanins  <= "0" & CLB_1_5_OUT_pin_2 & track_0_5_chanY_n0 & track_0_6_chanY_n1;
	track_1_5_chanX_n5_driver_mux_fanins  <= CLB_1_5_OUT_pin_2 & track_1_5_chanY_n2 & track_2_5_chanX_n5 & track_1_6_chanY_n13;
	track_1_5_chanX_n6_driver_mux_fanins  <= "0" & CLB_1_5_OUT_pin_2 & track_0_5_chanY_n2 & track_0_6_chanY_n3;
	track_1_5_chanX_n7_driver_mux_fanins  <= CLB_1_5_OUT_pin_2 & track_1_5_chanY_n4 & track_2_5_chanX_n7 & track_1_6_chanY_n11;
	track_1_5_chanX_n8_driver_mux_fanins  <= "0" & CLB_1_6_OUT_pin_0 & track_0_5_chanY_n4 & track_0_6_chanY_n5;
	track_1_5_chanX_n9_driver_mux_fanins  <= CLB_1_6_OUT_pin_0 & track_1_5_chanY_n6 & track_2_5_chanX_n9 & track_1_6_chanY_n9;
	track_1_5_chanY_n0_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_1_4_chanY_n0 & track_2_4_chanX_n3 & track_1_4_chanX_n0;
	track_1_5_chanY_n1_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_2_5_chanX_n13 & track_1_5_chanX_n2 & track_1_6_chanY_n1;
	track_1_5_chanY_n10_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_1_4_chanY_n10 & track_2_4_chanX_n13 & track_1_4_chanX_n6;
	track_1_5_chanY_n11_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_2_5_chanX_n3 & track_1_5_chanX_n12 & track_1_6_chanY_n11;
	track_1_5_chanY_n12_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_1_4_chanY_n12 & track_2_4_chanX_n15 & track_1_4_chanX_n4;
	track_1_5_chanY_n13_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_2_5_chanX_n1 & track_1_5_chanX_n14 & track_1_6_chanY_n13;
	track_1_5_chanY_n14_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_1_4_chanY_n14 & track_2_4_chanX_n1 & track_1_4_chanX_n2;
	track_1_5_chanY_n15_driver_mux_fanins <= CLB_2_5_OUT_pin_1 & track_2_5_chanX_n15 & track_1_5_chanX_n0 & track_1_6_chanY_n15;
	track_1_5_chanY_n2_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_1_4_chanY_n2 & track_2_4_chanX_n5 & track_1_4_chanX_n14;
	track_1_5_chanY_n3_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_2_5_chanX_n11 & track_1_5_chanX_n4 & track_1_6_chanY_n3;
	track_1_5_chanY_n4_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_1_4_chanY_n4 & track_2_4_chanX_n7 & track_1_4_chanX_n12;
	track_1_5_chanY_n5_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_2_5_chanX_n9 & track_1_5_chanX_n6 & track_1_6_chanY_n5;
	track_1_5_chanY_n6_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_1_4_chanY_n6 & track_2_4_chanX_n9 & track_1_4_chanX_n10;
	track_1_5_chanY_n7_driver_mux_fanins  <= CLB_1_5_OUT_pin_3 & track_2_5_chanX_n7 & track_1_5_chanX_n8 & track_1_6_chanY_n7;
	track_1_5_chanY_n8_driver_mux_fanins  <= CLB_2_5_OUT_pin_1 & track_1_4_chanY_n8 & track_2_4_chanX_n11 & track_1_4_chanX_n8;
	track_1_5_chanY_n9_driver_mux_fanins  <= CLB_2_5_OUT_pin_1 & track_2_5_chanX_n5 & track_1_5_chanX_n10 & track_1_6_chanY_n9;
	track_1_6_chanX_n0_driver_mux_fanins  <= "0" & IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_0_6_chanY_n12;
	track_1_6_chanX_n1_driver_mux_fanins  <= IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_1_6_chanY_n0 & track_2_6_chanX_n1;
	track_1_6_chanX_n10_driver_mux_fanins <= IO_1_7_OUT_pin_0 & track_0_6_chanY_n2;
	track_1_6_chanX_n11_driver_mux_fanins <= "0" & IO_1_7_OUT_pin_0 & track_1_6_chanY_n10 & track_2_6_chanX_n11;
	track_1_6_chanX_n12_driver_mux_fanins <= IO_1_7_OUT_pin_0 & track_0_6_chanY_n0;
	track_1_6_chanX_n13_driver_mux_fanins <= "0" & IO_1_7_OUT_pin_0 & track_1_6_chanY_n12 & track_2_6_chanX_n13;
	track_1_6_chanX_n14_driver_mux_fanins <= IO_1_7_OUT_pin_0 & track_0_6_chanY_n14;
	track_1_6_chanX_n15_driver_mux_fanins <= "0" & IO_1_7_OUT_pin_0 & track_1_6_chanY_n14 & track_2_6_chanX_n15;
	track_1_6_chanX_n2_driver_mux_fanins  <= "0" & IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_0_6_chanY_n10;
	track_1_6_chanX_n3_driver_mux_fanins  <= IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_1_6_chanY_n2 & track_2_6_chanX_n3;
	track_1_6_chanX_n4_driver_mux_fanins  <= "0" & IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_0_6_chanY_n8;
	track_1_6_chanX_n5_driver_mux_fanins  <= IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_1_6_chanY_n4 & track_2_6_chanX_n5;
	track_1_6_chanX_n6_driver_mux_fanins  <= "0" & IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_0_6_chanY_n6;
	track_1_6_chanX_n7_driver_mux_fanins  <= IO_1_7_OUT_pin_1 & CLB_1_6_OUT_pin_2 & track_1_6_chanY_n6 & track_2_6_chanX_n7;
	track_1_6_chanX_n8_driver_mux_fanins  <= IO_1_7_OUT_pin_0 & track_0_6_chanY_n4;
	track_1_6_chanX_n9_driver_mux_fanins  <= "0" & IO_1_7_OUT_pin_0 & track_1_6_chanY_n8 & track_2_6_chanX_n9;
	track_1_6_chanY_n0_driver_mux_fanins  <= CLB_1_6_OUT_pin_3 & track_1_5_chanY_n0 & track_2_5_chanX_n3 & track_1_5_chanX_n0;
	track_1_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_1_6_OUT_pin_3 & track_2_6_chanX_n1 & track_1_6_chanX_n0;
	track_1_6_chanY_n10_driver_mux_fanins <= CLB_2_6_OUT_pin_1 & track_1_5_chanY_n10 & track_2_5_chanX_n13 & track_1_5_chanX_n6;
	track_1_6_chanY_n11_driver_mux_fanins <= "0" & CLB_2_6_OUT_pin_1 & track_2_6_chanX_n5 & track_1_6_chanX_n4;
	track_1_6_chanY_n12_driver_mux_fanins <= CLB_2_6_OUT_pin_1 & track_1_5_chanY_n12 & track_2_5_chanX_n15 & track_1_5_chanX_n4;
	track_1_6_chanY_n13_driver_mux_fanins <= "0" & CLB_2_6_OUT_pin_1 & track_2_6_chanX_n7 & track_1_6_chanX_n6;
	track_1_6_chanY_n14_driver_mux_fanins <= CLB_2_6_OUT_pin_1 & track_1_5_chanY_n14 & track_2_5_chanX_n1 & track_1_5_chanX_n2;
	track_1_6_chanY_n15_driver_mux_fanins <= "0" & CLB_2_6_OUT_pin_1 & track_2_6_chanX_n15 & track_1_6_chanX_n14;
	track_1_6_chanY_n2_driver_mux_fanins  <= CLB_1_6_OUT_pin_3 & track_1_5_chanY_n2 & track_2_5_chanX_n5 & track_1_5_chanX_n14;
	track_1_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_1_6_OUT_pin_3 & track_2_6_chanX_n9 & track_1_6_chanX_n8;
	track_1_6_chanY_n4_driver_mux_fanins  <= CLB_1_6_OUT_pin_3 & track_1_5_chanY_n4 & track_2_5_chanX_n7 & track_1_5_chanX_n12;
	track_1_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_1_6_OUT_pin_3 & track_2_6_chanX_n11 & track_1_6_chanX_n10;
	track_1_6_chanY_n6_driver_mux_fanins  <= CLB_1_6_OUT_pin_3 & track_1_5_chanY_n6 & track_2_5_chanX_n9 & track_1_5_chanX_n10;
	track_1_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_1_6_OUT_pin_3 & track_2_6_chanX_n13 & track_1_6_chanX_n12;
	track_1_6_chanY_n8_driver_mux_fanins  <= CLB_2_6_OUT_pin_1 & track_1_5_chanY_n8 & track_2_5_chanX_n11 & track_1_5_chanX_n8;
	track_1_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_2_6_OUT_pin_1 & track_2_6_chanX_n3 & track_1_6_chanX_n2;
	track_2_0_chanX_n0_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_1_0_chanX_n0 & track_1_1_chanY_n1;
	track_2_0_chanX_n1_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_3_0_chanX_n1 & track_2_1_chanY_n1;
	track_2_0_chanX_n10_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_1_0_chanX_n10 & track_1_1_chanY_n11;
	track_2_0_chanX_n11_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_3_0_chanX_n11 & track_2_1_chanY_n11;
	track_2_0_chanX_n12_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_1_0_chanX_n12 & track_1_1_chanY_n13;
	track_2_0_chanX_n13_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_3_0_chanX_n13 & track_2_1_chanY_n13;
	track_2_0_chanX_n14_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_1_0_chanX_n14 & track_1_1_chanY_n15;
	track_2_0_chanX_n15_driver_mux_fanins <= "0" & IO_2_0_OUT_pin_1 & track_3_0_chanX_n15 & track_2_1_chanY_n15;
	track_2_0_chanX_n2_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_1_0_chanX_n2 & track_1_1_chanY_n3;
	track_2_0_chanX_n3_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_3_0_chanX_n3 & track_2_1_chanY_n3;
	track_2_0_chanX_n4_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_1_0_chanX_n4 & track_1_1_chanY_n5;
	track_2_0_chanX_n5_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_3_0_chanX_n5 & track_2_1_chanY_n5;
	track_2_0_chanX_n6_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_1_0_chanX_n6 & track_1_1_chanY_n7;
	track_2_0_chanX_n7_driver_mux_fanins  <= IO_2_0_OUT_pin_0 & CLB_2_1_OUT_pin_0 & track_3_0_chanX_n7 & track_2_1_chanY_n7;
	track_2_0_chanX_n8_driver_mux_fanins  <= "0" & IO_2_0_OUT_pin_1 & track_1_0_chanX_n8 & track_1_1_chanY_n9;
	track_2_0_chanX_n9_driver_mux_fanins  <= "0" & IO_2_0_OUT_pin_1 & track_3_0_chanX_n9 & track_2_1_chanY_n9;
	track_2_1_chanX_n0_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_1_1_chanY_n12 & track_1_1_chanX_n0 & track_1_2_chanY_n15;
	track_2_1_chanX_n1_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_2_1_chanY_n14 & track_3_1_chanX_n1 & track_2_2_chanY_n1;
	track_2_1_chanX_n10_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_1_1_chanY_n2 & track_1_1_chanX_n10 & track_1_2_chanY_n9;
	track_2_1_chanX_n11_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_2_1_chanY_n8 & track_3_1_chanX_n11 & track_2_2_chanY_n7;
	track_2_1_chanX_n12_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_1_1_chanY_n0 & track_1_1_chanX_n12 & track_1_2_chanY_n11;
	track_2_1_chanX_n13_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_2_1_chanY_n10 & track_3_1_chanX_n13 & track_2_2_chanY_n5;
	track_2_1_chanX_n14_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_1_1_chanY_n14 & track_1_1_chanX_n14 & track_1_2_chanY_n13;
	track_2_1_chanX_n15_driver_mux_fanins <= CLB_2_2_OUT_pin_0 & track_2_1_chanY_n12 & track_3_1_chanX_n15 & track_2_2_chanY_n3;
	track_2_1_chanX_n2_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_1_1_chanY_n10 & track_1_1_chanX_n2 & track_1_2_chanY_n1;
	track_2_1_chanX_n3_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_2_1_chanY_n0 & track_3_1_chanX_n3 & track_2_2_chanY_n15;
	track_2_1_chanX_n4_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_1_1_chanY_n8 & track_1_1_chanX_n4 & track_1_2_chanY_n3;
	track_2_1_chanX_n5_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_2_1_chanY_n2 & track_3_1_chanX_n5 & track_2_2_chanY_n13;
	track_2_1_chanX_n6_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_1_1_chanY_n6 & track_1_1_chanX_n6 & track_1_2_chanY_n5;
	track_2_1_chanX_n7_driver_mux_fanins  <= CLB_2_1_OUT_pin_2 & track_2_1_chanY_n4 & track_3_1_chanX_n7 & track_2_2_chanY_n11;
	track_2_1_chanX_n8_driver_mux_fanins  <= CLB_2_2_OUT_pin_0 & track_1_1_chanY_n4 & track_1_1_chanX_n8 & track_1_2_chanY_n7;
	track_2_1_chanX_n9_driver_mux_fanins  <= CLB_2_2_OUT_pin_0 & track_2_1_chanY_n6 & track_3_1_chanX_n9 & track_2_2_chanY_n9;
	track_2_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_2_1_OUT_pin_3 & track_3_0_chanX_n7 & track_2_0_chanX_n6;
	track_2_1_chanY_n1_driver_mux_fanins  <= CLB_2_1_OUT_pin_3 & track_3_1_chanX_n13 & track_2_1_chanX_n2 & track_2_2_chanY_n1;
	track_2_1_chanY_n10_driver_mux_fanins <= "0" & CLB_3_1_OUT_pin_1 & track_3_0_chanX_n11 & track_2_0_chanX_n10;
	track_2_1_chanY_n11_driver_mux_fanins <= CLB_3_1_OUT_pin_1 & track_3_1_chanX_n3 & track_2_1_chanX_n12 & track_2_2_chanY_n11;
	track_2_1_chanY_n12_driver_mux_fanins <= "0" & CLB_3_1_OUT_pin_1 & track_3_0_chanX_n13 & track_2_0_chanX_n12;
	track_2_1_chanY_n13_driver_mux_fanins <= CLB_3_1_OUT_pin_1 & track_3_1_chanX_n1 & track_2_1_chanX_n14 & track_2_2_chanY_n13;
	track_2_1_chanY_n14_driver_mux_fanins <= "0" & CLB_3_1_OUT_pin_1 & track_3_0_chanX_n15 & track_2_0_chanX_n14;
	track_2_1_chanY_n15_driver_mux_fanins <= CLB_3_1_OUT_pin_1 & track_3_1_chanX_n15 & track_2_1_chanX_n0 & track_2_2_chanY_n15;
	track_2_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_2_1_OUT_pin_3 & track_3_0_chanX_n9 & track_2_0_chanX_n8;
	track_2_1_chanY_n3_driver_mux_fanins  <= CLB_2_1_OUT_pin_3 & track_3_1_chanX_n11 & track_2_1_chanX_n4 & track_2_2_chanY_n3;
	track_2_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_2_1_OUT_pin_3 & track_3_0_chanX_n1 & track_2_0_chanX_n0;
	track_2_1_chanY_n5_driver_mux_fanins  <= CLB_2_1_OUT_pin_3 & track_3_1_chanX_n9 & track_2_1_chanX_n6 & track_2_2_chanY_n5;
	track_2_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_2_1_OUT_pin_3 & track_3_0_chanX_n3 & track_2_0_chanX_n2;
	track_2_1_chanY_n7_driver_mux_fanins  <= CLB_2_1_OUT_pin_3 & track_3_1_chanX_n7 & track_2_1_chanX_n8 & track_2_2_chanY_n7;
	track_2_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_3_1_OUT_pin_1 & track_3_0_chanX_n5 & track_2_0_chanX_n4;
	track_2_1_chanY_n9_driver_mux_fanins  <= CLB_3_1_OUT_pin_1 & track_3_1_chanX_n5 & track_2_1_chanX_n10 & track_2_2_chanY_n9;
	track_2_2_chanX_n0_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_1_2_chanY_n12 & track_1_2_chanX_n0 & track_1_3_chanY_n15;
	track_2_2_chanX_n1_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_2_2_chanY_n14 & track_3_2_chanX_n1 & track_2_3_chanY_n1;
	track_2_2_chanX_n10_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_1_2_chanY_n2 & track_1_2_chanX_n10 & track_1_3_chanY_n9;
	track_2_2_chanX_n11_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_2_2_chanY_n8 & track_3_2_chanX_n11 & track_2_3_chanY_n7;
	track_2_2_chanX_n12_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_1_2_chanY_n0 & track_1_2_chanX_n12 & track_1_3_chanY_n11;
	track_2_2_chanX_n13_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_2_2_chanY_n10 & track_3_2_chanX_n13 & track_2_3_chanY_n5;
	track_2_2_chanX_n14_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_1_2_chanY_n14 & track_1_2_chanX_n14 & track_1_3_chanY_n13;
	track_2_2_chanX_n15_driver_mux_fanins <= CLB_2_3_OUT_pin_0 & track_2_2_chanY_n12 & track_3_2_chanX_n15 & track_2_3_chanY_n3;
	track_2_2_chanX_n2_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_1_2_chanY_n10 & track_1_2_chanX_n2 & track_1_3_chanY_n1;
	track_2_2_chanX_n3_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_2_2_chanY_n0 & track_3_2_chanX_n3 & track_2_3_chanY_n15;
	track_2_2_chanX_n4_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_1_2_chanY_n8 & track_1_2_chanX_n4 & track_1_3_chanY_n3;
	track_2_2_chanX_n5_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_2_2_chanY_n2 & track_3_2_chanX_n5 & track_2_3_chanY_n13;
	track_2_2_chanX_n6_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_1_2_chanY_n6 & track_1_2_chanX_n6 & track_1_3_chanY_n5;
	track_2_2_chanX_n7_driver_mux_fanins  <= CLB_2_2_OUT_pin_2 & track_2_2_chanY_n4 & track_3_2_chanX_n7 & track_2_3_chanY_n11;
	track_2_2_chanX_n8_driver_mux_fanins  <= CLB_2_3_OUT_pin_0 & track_1_2_chanY_n4 & track_1_2_chanX_n8 & track_1_3_chanY_n7;
	track_2_2_chanX_n9_driver_mux_fanins  <= CLB_2_3_OUT_pin_0 & track_2_2_chanY_n6 & track_3_2_chanX_n9 & track_2_3_chanY_n9;
	track_2_2_chanY_n0_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_2_1_chanY_n0 & track_3_1_chanX_n3 & track_2_1_chanX_n0;
	track_2_2_chanY_n1_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_3_2_chanX_n13 & track_2_2_chanX_n2 & track_2_3_chanY_n1;
	track_2_2_chanY_n10_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_2_1_chanY_n10 & track_3_1_chanX_n13 & track_2_1_chanX_n6;
	track_2_2_chanY_n11_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_3_2_chanX_n3 & track_2_2_chanX_n12 & track_2_3_chanY_n11;
	track_2_2_chanY_n12_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_2_1_chanY_n12 & track_3_1_chanX_n15 & track_2_1_chanX_n4;
	track_2_2_chanY_n13_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_3_2_chanX_n1 & track_2_2_chanX_n14 & track_2_3_chanY_n13;
	track_2_2_chanY_n14_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_2_1_chanY_n14 & track_3_1_chanX_n1 & track_2_1_chanX_n2;
	track_2_2_chanY_n15_driver_mux_fanins <= CLB_3_2_OUT_pin_1 & track_3_2_chanX_n15 & track_2_2_chanX_n0 & track_2_3_chanY_n15;
	track_2_2_chanY_n2_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_2_1_chanY_n2 & track_3_1_chanX_n5 & track_2_1_chanX_n14;
	track_2_2_chanY_n3_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_3_2_chanX_n11 & track_2_2_chanX_n4 & track_2_3_chanY_n3;
	track_2_2_chanY_n4_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_2_1_chanY_n4 & track_3_1_chanX_n7 & track_2_1_chanX_n12;
	track_2_2_chanY_n5_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_3_2_chanX_n9 & track_2_2_chanX_n6 & track_2_3_chanY_n5;
	track_2_2_chanY_n6_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_2_1_chanY_n6 & track_3_1_chanX_n9 & track_2_1_chanX_n10;
	track_2_2_chanY_n7_driver_mux_fanins  <= CLB_2_2_OUT_pin_3 & track_3_2_chanX_n7 & track_2_2_chanX_n8 & track_2_3_chanY_n7;
	track_2_2_chanY_n8_driver_mux_fanins  <= CLB_3_2_OUT_pin_1 & track_2_1_chanY_n8 & track_3_1_chanX_n11 & track_2_1_chanX_n8;
	track_2_2_chanY_n9_driver_mux_fanins  <= CLB_3_2_OUT_pin_1 & track_3_2_chanX_n5 & track_2_2_chanX_n10 & track_2_3_chanY_n9;
	track_2_3_chanX_n0_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_1_3_chanY_n12 & track_1_3_chanX_n0 & track_1_4_chanY_n15;
	track_2_3_chanX_n1_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_2_3_chanY_n14 & track_3_3_chanX_n1 & track_2_4_chanY_n1;
	track_2_3_chanX_n10_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_1_3_chanY_n2 & track_1_3_chanX_n10 & track_1_4_chanY_n9;
	track_2_3_chanX_n11_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_2_3_chanY_n8 & track_3_3_chanX_n11 & track_2_4_chanY_n7;
	track_2_3_chanX_n12_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_1_3_chanY_n0 & track_1_3_chanX_n12 & track_1_4_chanY_n11;
	track_2_3_chanX_n13_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_2_3_chanY_n10 & track_3_3_chanX_n13 & track_2_4_chanY_n5;
	track_2_3_chanX_n14_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_1_3_chanY_n14 & track_1_3_chanX_n14 & track_1_4_chanY_n13;
	track_2_3_chanX_n15_driver_mux_fanins <= CLB_2_4_OUT_pin_0 & track_2_3_chanY_n12 & track_3_3_chanX_n15 & track_2_4_chanY_n3;
	track_2_3_chanX_n2_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_1_3_chanY_n10 & track_1_3_chanX_n2 & track_1_4_chanY_n1;
	track_2_3_chanX_n3_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_2_3_chanY_n0 & track_3_3_chanX_n3 & track_2_4_chanY_n15;
	track_2_3_chanX_n4_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_1_3_chanY_n8 & track_1_3_chanX_n4 & track_1_4_chanY_n3;
	track_2_3_chanX_n5_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_2_3_chanY_n2 & track_3_3_chanX_n5 & track_2_4_chanY_n13;
	track_2_3_chanX_n6_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_1_3_chanY_n6 & track_1_3_chanX_n6 & track_1_4_chanY_n5;
	track_2_3_chanX_n7_driver_mux_fanins  <= CLB_2_3_OUT_pin_2 & track_2_3_chanY_n4 & track_3_3_chanX_n7 & track_2_4_chanY_n11;
	track_2_3_chanX_n8_driver_mux_fanins  <= CLB_2_4_OUT_pin_0 & track_1_3_chanY_n4 & track_1_3_chanX_n8 & track_1_4_chanY_n7;
	track_2_3_chanX_n9_driver_mux_fanins  <= CLB_2_4_OUT_pin_0 & track_2_3_chanY_n6 & track_3_3_chanX_n9 & track_2_4_chanY_n9;
	track_2_3_chanY_n0_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_2_2_chanY_n0 & track_3_2_chanX_n3 & track_2_2_chanX_n0;
	track_2_3_chanY_n1_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_3_3_chanX_n13 & track_2_3_chanX_n2 & track_2_4_chanY_n1;
	track_2_3_chanY_n10_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_2_2_chanY_n10 & track_3_2_chanX_n13 & track_2_2_chanX_n6;
	track_2_3_chanY_n11_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_3_3_chanX_n3 & track_2_3_chanX_n12 & track_2_4_chanY_n11;
	track_2_3_chanY_n12_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_2_2_chanY_n12 & track_3_2_chanX_n15 & track_2_2_chanX_n4;
	track_2_3_chanY_n13_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_3_3_chanX_n1 & track_2_3_chanX_n14 & track_2_4_chanY_n13;
	track_2_3_chanY_n14_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_2_2_chanY_n14 & track_3_2_chanX_n1 & track_2_2_chanX_n2;
	track_2_3_chanY_n15_driver_mux_fanins <= CLB_3_3_OUT_pin_1 & track_3_3_chanX_n15 & track_2_3_chanX_n0 & track_2_4_chanY_n15;
	track_2_3_chanY_n2_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_2_2_chanY_n2 & track_3_2_chanX_n5 & track_2_2_chanX_n14;
	track_2_3_chanY_n3_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_3_3_chanX_n11 & track_2_3_chanX_n4 & track_2_4_chanY_n3;
	track_2_3_chanY_n4_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_2_2_chanY_n4 & track_3_2_chanX_n7 & track_2_2_chanX_n12;
	track_2_3_chanY_n5_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_3_3_chanX_n9 & track_2_3_chanX_n6 & track_2_4_chanY_n5;
	track_2_3_chanY_n6_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_2_2_chanY_n6 & track_3_2_chanX_n9 & track_2_2_chanX_n10;
	track_2_3_chanY_n7_driver_mux_fanins  <= CLB_2_3_OUT_pin_3 & track_3_3_chanX_n7 & track_2_3_chanX_n8 & track_2_4_chanY_n7;
	track_2_3_chanY_n8_driver_mux_fanins  <= CLB_3_3_OUT_pin_1 & track_2_2_chanY_n8 & track_3_2_chanX_n11 & track_2_2_chanX_n8;
	track_2_3_chanY_n9_driver_mux_fanins  <= CLB_3_3_OUT_pin_1 & track_3_3_chanX_n5 & track_2_3_chanX_n10 & track_2_4_chanY_n9;
	track_2_4_chanX_n0_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_1_4_chanY_n12 & track_1_4_chanX_n0 & track_1_5_chanY_n15;
	track_2_4_chanX_n1_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_2_4_chanY_n14 & track_3_4_chanX_n1 & track_2_5_chanY_n1;
	track_2_4_chanX_n10_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_1_4_chanY_n2 & track_1_4_chanX_n10 & track_1_5_chanY_n9;
	track_2_4_chanX_n11_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_2_4_chanY_n8 & track_3_4_chanX_n11 & track_2_5_chanY_n7;
	track_2_4_chanX_n12_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_1_4_chanY_n0 & track_1_4_chanX_n12 & track_1_5_chanY_n11;
	track_2_4_chanX_n13_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_2_4_chanY_n10 & track_3_4_chanX_n13 & track_2_5_chanY_n5;
	track_2_4_chanX_n14_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_1_4_chanY_n14 & track_1_4_chanX_n14 & track_1_5_chanY_n13;
	track_2_4_chanX_n15_driver_mux_fanins <= CLB_2_5_OUT_pin_0 & track_2_4_chanY_n12 & track_3_4_chanX_n15 & track_2_5_chanY_n3;
	track_2_4_chanX_n2_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_1_4_chanY_n10 & track_1_4_chanX_n2 & track_1_5_chanY_n1;
	track_2_4_chanX_n3_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_2_4_chanY_n0 & track_3_4_chanX_n3 & track_2_5_chanY_n15;
	track_2_4_chanX_n4_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_1_4_chanY_n8 & track_1_4_chanX_n4 & track_1_5_chanY_n3;
	track_2_4_chanX_n5_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_2_4_chanY_n2 & track_3_4_chanX_n5 & track_2_5_chanY_n13;
	track_2_4_chanX_n6_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_1_4_chanY_n6 & track_1_4_chanX_n6 & track_1_5_chanY_n5;
	track_2_4_chanX_n7_driver_mux_fanins  <= CLB_2_4_OUT_pin_2 & track_2_4_chanY_n4 & track_3_4_chanX_n7 & track_2_5_chanY_n11;
	track_2_4_chanX_n8_driver_mux_fanins  <= CLB_2_5_OUT_pin_0 & track_1_4_chanY_n4 & track_1_4_chanX_n8 & track_1_5_chanY_n7;
	track_2_4_chanX_n9_driver_mux_fanins  <= CLB_2_5_OUT_pin_0 & track_2_4_chanY_n6 & track_3_4_chanX_n9 & track_2_5_chanY_n9;
	track_2_4_chanY_n0_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_2_3_chanY_n0 & track_3_3_chanX_n3 & track_2_3_chanX_n0;
	track_2_4_chanY_n1_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_3_4_chanX_n13 & track_2_4_chanX_n2 & track_2_5_chanY_n1;
	track_2_4_chanY_n10_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_2_3_chanY_n10 & track_3_3_chanX_n13 & track_2_3_chanX_n6;
	track_2_4_chanY_n11_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_3_4_chanX_n3 & track_2_4_chanX_n12 & track_2_5_chanY_n11;
	track_2_4_chanY_n12_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_2_3_chanY_n12 & track_3_3_chanX_n15 & track_2_3_chanX_n4;
	track_2_4_chanY_n13_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_3_4_chanX_n1 & track_2_4_chanX_n14 & track_2_5_chanY_n13;
	track_2_4_chanY_n14_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_2_3_chanY_n14 & track_3_3_chanX_n1 & track_2_3_chanX_n2;
	track_2_4_chanY_n15_driver_mux_fanins <= CLB_3_4_OUT_pin_1 & track_3_4_chanX_n15 & track_2_4_chanX_n0 & track_2_5_chanY_n15;
	track_2_4_chanY_n2_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_2_3_chanY_n2 & track_3_3_chanX_n5 & track_2_3_chanX_n14;
	track_2_4_chanY_n3_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_3_4_chanX_n11 & track_2_4_chanX_n4 & track_2_5_chanY_n3;
	track_2_4_chanY_n4_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_2_3_chanY_n4 & track_3_3_chanX_n7 & track_2_3_chanX_n12;
	track_2_4_chanY_n5_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_3_4_chanX_n9 & track_2_4_chanX_n6 & track_2_5_chanY_n5;
	track_2_4_chanY_n6_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_2_3_chanY_n6 & track_3_3_chanX_n9 & track_2_3_chanX_n10;
	track_2_4_chanY_n7_driver_mux_fanins  <= CLB_2_4_OUT_pin_3 & track_3_4_chanX_n7 & track_2_4_chanX_n8 & track_2_5_chanY_n7;
	track_2_4_chanY_n8_driver_mux_fanins  <= CLB_3_4_OUT_pin_1 & track_2_3_chanY_n8 & track_3_3_chanX_n11 & track_2_3_chanX_n8;
	track_2_4_chanY_n9_driver_mux_fanins  <= CLB_3_4_OUT_pin_1 & track_3_4_chanX_n5 & track_2_4_chanX_n10 & track_2_5_chanY_n9;
	track_2_5_chanX_n0_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_1_5_chanY_n12 & track_1_5_chanX_n0 & track_1_6_chanY_n15;
	track_2_5_chanX_n1_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_2_5_chanY_n14 & track_3_5_chanX_n1 & track_2_6_chanY_n1;
	track_2_5_chanX_n10_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_1_5_chanY_n2 & track_1_5_chanX_n10 & track_1_6_chanY_n9;
	track_2_5_chanX_n11_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_2_5_chanY_n8 & track_3_5_chanX_n11 & track_2_6_chanY_n7;
	track_2_5_chanX_n12_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_1_5_chanY_n0 & track_1_5_chanX_n12 & track_1_6_chanY_n11;
	track_2_5_chanX_n13_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_2_5_chanY_n10 & track_3_5_chanX_n13 & track_2_6_chanY_n5;
	track_2_5_chanX_n14_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_1_5_chanY_n14 & track_1_5_chanX_n14 & track_1_6_chanY_n13;
	track_2_5_chanX_n15_driver_mux_fanins <= CLB_2_6_OUT_pin_0 & track_2_5_chanY_n12 & track_3_5_chanX_n15 & track_2_6_chanY_n3;
	track_2_5_chanX_n2_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_1_5_chanY_n10 & track_1_5_chanX_n2 & track_1_6_chanY_n1;
	track_2_5_chanX_n3_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_2_5_chanY_n0 & track_3_5_chanX_n3 & track_2_6_chanY_n15;
	track_2_5_chanX_n4_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_1_5_chanY_n8 & track_1_5_chanX_n4 & track_1_6_chanY_n3;
	track_2_5_chanX_n5_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_2_5_chanY_n2 & track_3_5_chanX_n5 & track_2_6_chanY_n13;
	track_2_5_chanX_n6_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_1_5_chanY_n6 & track_1_5_chanX_n6 & track_1_6_chanY_n5;
	track_2_5_chanX_n7_driver_mux_fanins  <= CLB_2_5_OUT_pin_2 & track_2_5_chanY_n4 & track_3_5_chanX_n7 & track_2_6_chanY_n11;
	track_2_5_chanX_n8_driver_mux_fanins  <= CLB_2_6_OUT_pin_0 & track_1_5_chanY_n4 & track_1_5_chanX_n8 & track_1_6_chanY_n7;
	track_2_5_chanX_n9_driver_mux_fanins  <= CLB_2_6_OUT_pin_0 & track_2_5_chanY_n6 & track_3_5_chanX_n9 & track_2_6_chanY_n9;
	track_2_5_chanY_n0_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_2_4_chanY_n0 & track_3_4_chanX_n3 & track_2_4_chanX_n0;
	track_2_5_chanY_n1_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_3_5_chanX_n13 & track_2_5_chanX_n2 & track_2_6_chanY_n1;
	track_2_5_chanY_n10_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_2_4_chanY_n10 & track_3_4_chanX_n13 & track_2_4_chanX_n6;
	track_2_5_chanY_n11_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_3_5_chanX_n3 & track_2_5_chanX_n12 & track_2_6_chanY_n11;
	track_2_5_chanY_n12_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_2_4_chanY_n12 & track_3_4_chanX_n15 & track_2_4_chanX_n4;
	track_2_5_chanY_n13_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_3_5_chanX_n1 & track_2_5_chanX_n14 & track_2_6_chanY_n13;
	track_2_5_chanY_n14_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_2_4_chanY_n14 & track_3_4_chanX_n1 & track_2_4_chanX_n2;
	track_2_5_chanY_n15_driver_mux_fanins <= CLB_3_5_OUT_pin_1 & track_3_5_chanX_n15 & track_2_5_chanX_n0 & track_2_6_chanY_n15;
	track_2_5_chanY_n2_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_2_4_chanY_n2 & track_3_4_chanX_n5 & track_2_4_chanX_n14;
	track_2_5_chanY_n3_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_3_5_chanX_n11 & track_2_5_chanX_n4 & track_2_6_chanY_n3;
	track_2_5_chanY_n4_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_2_4_chanY_n4 & track_3_4_chanX_n7 & track_2_4_chanX_n12;
	track_2_5_chanY_n5_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_3_5_chanX_n9 & track_2_5_chanX_n6 & track_2_6_chanY_n5;
	track_2_5_chanY_n6_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_2_4_chanY_n6 & track_3_4_chanX_n9 & track_2_4_chanX_n10;
	track_2_5_chanY_n7_driver_mux_fanins  <= CLB_2_5_OUT_pin_3 & track_3_5_chanX_n7 & track_2_5_chanX_n8 & track_2_6_chanY_n7;
	track_2_5_chanY_n8_driver_mux_fanins  <= CLB_3_5_OUT_pin_1 & track_2_4_chanY_n8 & track_3_4_chanX_n11 & track_2_4_chanX_n8;
	track_2_5_chanY_n9_driver_mux_fanins  <= CLB_3_5_OUT_pin_1 & track_3_5_chanX_n5 & track_2_5_chanX_n10 & track_2_6_chanY_n9;
	track_2_6_chanX_n0_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_1_6_chanY_n0 & track_1_6_chanX_n0;
	track_2_6_chanX_n1_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_2_6_chanY_n0 & track_3_6_chanX_n1;
	track_2_6_chanX_n10_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_1_6_chanY_n10 & track_1_6_chanX_n10;
	track_2_6_chanX_n11_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_2_6_chanY_n10 & track_3_6_chanX_n11;
	track_2_6_chanX_n12_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_1_6_chanY_n12 & track_1_6_chanX_n12;
	track_2_6_chanX_n13_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_2_6_chanY_n12 & track_3_6_chanX_n13;
	track_2_6_chanX_n14_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_1_6_chanY_n14 & track_1_6_chanX_n14;
	track_2_6_chanX_n15_driver_mux_fanins <= "0" & IO_2_7_OUT_pin_0 & track_2_6_chanY_n14 & track_3_6_chanX_n15;
	track_2_6_chanX_n2_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_1_6_chanY_n2 & track_1_6_chanX_n2;
	track_2_6_chanX_n3_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_2_6_chanY_n2 & track_3_6_chanX_n3;
	track_2_6_chanX_n4_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_1_6_chanY_n4 & track_1_6_chanX_n4;
	track_2_6_chanX_n5_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_2_6_chanY_n4 & track_3_6_chanX_n5;
	track_2_6_chanX_n6_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_1_6_chanY_n6 & track_1_6_chanX_n6;
	track_2_6_chanX_n7_driver_mux_fanins  <= IO_2_7_OUT_pin_1 & CLB_2_6_OUT_pin_2 & track_2_6_chanY_n6 & track_3_6_chanX_n7;
	track_2_6_chanX_n8_driver_mux_fanins  <= "0" & IO_2_7_OUT_pin_0 & track_1_6_chanY_n8 & track_1_6_chanX_n8;
	track_2_6_chanX_n9_driver_mux_fanins  <= "0" & IO_2_7_OUT_pin_0 & track_2_6_chanY_n8 & track_3_6_chanX_n9;
	track_2_6_chanY_n0_driver_mux_fanins  <= CLB_2_6_OUT_pin_3 & track_2_5_chanY_n0 & track_3_5_chanX_n3 & track_2_5_chanX_n0;
	track_2_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_2_6_OUT_pin_3 & track_3_6_chanX_n1 & track_2_6_chanX_n0;
	track_2_6_chanY_n10_driver_mux_fanins <= CLB_3_6_OUT_pin_1 & track_2_5_chanY_n10 & track_3_5_chanX_n13 & track_2_5_chanX_n6;
	track_2_6_chanY_n11_driver_mux_fanins <= "0" & CLB_3_6_OUT_pin_1 & track_3_6_chanX_n5 & track_2_6_chanX_n4;
	track_2_6_chanY_n12_driver_mux_fanins <= CLB_3_6_OUT_pin_1 & track_2_5_chanY_n12 & track_3_5_chanX_n15 & track_2_5_chanX_n4;
	track_2_6_chanY_n13_driver_mux_fanins <= "0" & CLB_3_6_OUT_pin_1 & track_3_6_chanX_n7 & track_2_6_chanX_n6;
	track_2_6_chanY_n14_driver_mux_fanins <= CLB_3_6_OUT_pin_1 & track_2_5_chanY_n14 & track_3_5_chanX_n1 & track_2_5_chanX_n2;
	track_2_6_chanY_n15_driver_mux_fanins <= "0" & CLB_3_6_OUT_pin_1 & track_3_6_chanX_n15 & track_2_6_chanX_n14;
	track_2_6_chanY_n2_driver_mux_fanins  <= CLB_2_6_OUT_pin_3 & track_2_5_chanY_n2 & track_3_5_chanX_n5 & track_2_5_chanX_n14;
	track_2_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_2_6_OUT_pin_3 & track_3_6_chanX_n9 & track_2_6_chanX_n8;
	track_2_6_chanY_n4_driver_mux_fanins  <= CLB_2_6_OUT_pin_3 & track_2_5_chanY_n4 & track_3_5_chanX_n7 & track_2_5_chanX_n12;
	track_2_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_2_6_OUT_pin_3 & track_3_6_chanX_n11 & track_2_6_chanX_n10;
	track_2_6_chanY_n6_driver_mux_fanins  <= CLB_2_6_OUT_pin_3 & track_2_5_chanY_n6 & track_3_5_chanX_n9 & track_2_5_chanX_n10;
	track_2_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_2_6_OUT_pin_3 & track_3_6_chanX_n13 & track_2_6_chanX_n12;
	track_2_6_chanY_n8_driver_mux_fanins  <= CLB_3_6_OUT_pin_1 & track_2_5_chanY_n8 & track_3_5_chanX_n11 & track_2_5_chanX_n8;
	track_2_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_3_6_OUT_pin_1 & track_3_6_chanX_n3 & track_2_6_chanX_n2;
	track_3_0_chanX_n0_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_2_0_chanX_n0 & track_2_1_chanY_n1;
	track_3_0_chanX_n1_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_4_0_chanX_n1 & track_3_1_chanY_n1;
	track_3_0_chanX_n10_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_2_0_chanX_n10 & track_2_1_chanY_n11;
	track_3_0_chanX_n11_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_4_0_chanX_n11 & track_3_1_chanY_n11;
	track_3_0_chanX_n12_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_2_0_chanX_n12 & track_2_1_chanY_n13;
	track_3_0_chanX_n13_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_4_0_chanX_n13 & track_3_1_chanY_n13;
	track_3_0_chanX_n14_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_2_0_chanX_n14 & track_2_1_chanY_n15;
	track_3_0_chanX_n15_driver_mux_fanins <= "0" & IO_3_0_OUT_pin_1 & track_4_0_chanX_n15 & track_3_1_chanY_n15;
	track_3_0_chanX_n2_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_2_0_chanX_n2 & track_2_1_chanY_n3;
	track_3_0_chanX_n3_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_4_0_chanX_n3 & track_3_1_chanY_n3;
	track_3_0_chanX_n4_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_2_0_chanX_n4 & track_2_1_chanY_n5;
	track_3_0_chanX_n5_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_4_0_chanX_n5 & track_3_1_chanY_n5;
	track_3_0_chanX_n6_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_2_0_chanX_n6 & track_2_1_chanY_n7;
	track_3_0_chanX_n7_driver_mux_fanins  <= IO_3_0_OUT_pin_0 & CLB_3_1_OUT_pin_0 & track_4_0_chanX_n7 & track_3_1_chanY_n7;
	track_3_0_chanX_n8_driver_mux_fanins  <= "0" & IO_3_0_OUT_pin_1 & track_2_0_chanX_n8 & track_2_1_chanY_n9;
	track_3_0_chanX_n9_driver_mux_fanins  <= "0" & IO_3_0_OUT_pin_1 & track_4_0_chanX_n9 & track_3_1_chanY_n9;
	track_3_1_chanX_n0_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_2_1_chanY_n12 & track_2_1_chanX_n0 & track_2_2_chanY_n15;
	track_3_1_chanX_n1_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_3_1_chanY_n14 & track_4_1_chanX_n1 & track_3_2_chanY_n1;
	track_3_1_chanX_n10_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_2_1_chanY_n2 & track_2_1_chanX_n10 & track_2_2_chanY_n9;
	track_3_1_chanX_n11_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_3_1_chanY_n8 & track_4_1_chanX_n11 & track_3_2_chanY_n7;
	track_3_1_chanX_n12_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_2_1_chanY_n0 & track_2_1_chanX_n12 & track_2_2_chanY_n11;
	track_3_1_chanX_n13_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_3_1_chanY_n10 & track_4_1_chanX_n13 & track_3_2_chanY_n5;
	track_3_1_chanX_n14_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_2_1_chanY_n14 & track_2_1_chanX_n14 & track_2_2_chanY_n13;
	track_3_1_chanX_n15_driver_mux_fanins <= CLB_3_2_OUT_pin_0 & track_3_1_chanY_n12 & track_4_1_chanX_n15 & track_3_2_chanY_n3;
	track_3_1_chanX_n2_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_2_1_chanY_n10 & track_2_1_chanX_n2 & track_2_2_chanY_n1;
	track_3_1_chanX_n3_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_3_1_chanY_n0 & track_4_1_chanX_n3 & track_3_2_chanY_n15;
	track_3_1_chanX_n4_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_2_1_chanY_n8 & track_2_1_chanX_n4 & track_2_2_chanY_n3;
	track_3_1_chanX_n5_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_3_1_chanY_n2 & track_4_1_chanX_n5 & track_3_2_chanY_n13;
	track_3_1_chanX_n6_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_2_1_chanY_n6 & track_2_1_chanX_n6 & track_2_2_chanY_n5;
	track_3_1_chanX_n7_driver_mux_fanins  <= CLB_3_1_OUT_pin_2 & track_3_1_chanY_n4 & track_4_1_chanX_n7 & track_3_2_chanY_n11;
	track_3_1_chanX_n8_driver_mux_fanins  <= CLB_3_2_OUT_pin_0 & track_2_1_chanY_n4 & track_2_1_chanX_n8 & track_2_2_chanY_n7;
	track_3_1_chanX_n9_driver_mux_fanins  <= CLB_3_2_OUT_pin_0 & track_3_1_chanY_n6 & track_4_1_chanX_n9 & track_3_2_chanY_n9;
	track_3_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_3_1_OUT_pin_3 & track_4_0_chanX_n7 & track_3_0_chanX_n6;
	track_3_1_chanY_n1_driver_mux_fanins  <= CLB_3_1_OUT_pin_3 & track_4_1_chanX_n13 & track_3_1_chanX_n2 & track_3_2_chanY_n1;
	track_3_1_chanY_n10_driver_mux_fanins <= "0" & CLB_4_1_OUT_pin_1 & track_4_0_chanX_n11 & track_3_0_chanX_n10;
	track_3_1_chanY_n11_driver_mux_fanins <= CLB_4_1_OUT_pin_1 & track_4_1_chanX_n3 & track_3_1_chanX_n12 & track_3_2_chanY_n11;
	track_3_1_chanY_n12_driver_mux_fanins <= "0" & CLB_4_1_OUT_pin_1 & track_4_0_chanX_n13 & track_3_0_chanX_n12;
	track_3_1_chanY_n13_driver_mux_fanins <= CLB_4_1_OUT_pin_1 & track_4_1_chanX_n1 & track_3_1_chanX_n14 & track_3_2_chanY_n13;
	track_3_1_chanY_n14_driver_mux_fanins <= "0" & CLB_4_1_OUT_pin_1 & track_4_0_chanX_n15 & track_3_0_chanX_n14;
	track_3_1_chanY_n15_driver_mux_fanins <= CLB_4_1_OUT_pin_1 & track_4_1_chanX_n15 & track_3_1_chanX_n0 & track_3_2_chanY_n15;
	track_3_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_3_1_OUT_pin_3 & track_4_0_chanX_n9 & track_3_0_chanX_n8;
	track_3_1_chanY_n3_driver_mux_fanins  <= CLB_3_1_OUT_pin_3 & track_4_1_chanX_n11 & track_3_1_chanX_n4 & track_3_2_chanY_n3;
	track_3_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_3_1_OUT_pin_3 & track_4_0_chanX_n1 & track_3_0_chanX_n0;
	track_3_1_chanY_n5_driver_mux_fanins  <= CLB_3_1_OUT_pin_3 & track_4_1_chanX_n9 & track_3_1_chanX_n6 & track_3_2_chanY_n5;
	track_3_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_3_1_OUT_pin_3 & track_4_0_chanX_n3 & track_3_0_chanX_n2;
	track_3_1_chanY_n7_driver_mux_fanins  <= CLB_3_1_OUT_pin_3 & track_4_1_chanX_n7 & track_3_1_chanX_n8 & track_3_2_chanY_n7;
	track_3_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_4_1_OUT_pin_1 & track_4_0_chanX_n5 & track_3_0_chanX_n4;
	track_3_1_chanY_n9_driver_mux_fanins  <= CLB_4_1_OUT_pin_1 & track_4_1_chanX_n5 & track_3_1_chanX_n10 & track_3_2_chanY_n9;
	track_3_2_chanX_n0_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_2_2_chanY_n12 & track_2_2_chanX_n0 & track_2_3_chanY_n15;
	track_3_2_chanX_n1_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_3_2_chanY_n14 & track_4_2_chanX_n1 & track_3_3_chanY_n1;
	track_3_2_chanX_n10_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_2_2_chanY_n2 & track_2_2_chanX_n10 & track_2_3_chanY_n9;
	track_3_2_chanX_n11_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_3_2_chanY_n8 & track_4_2_chanX_n11 & track_3_3_chanY_n7;
	track_3_2_chanX_n12_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_2_2_chanY_n0 & track_2_2_chanX_n12 & track_2_3_chanY_n11;
	track_3_2_chanX_n13_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_3_2_chanY_n10 & track_4_2_chanX_n13 & track_3_3_chanY_n5;
	track_3_2_chanX_n14_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_2_2_chanY_n14 & track_2_2_chanX_n14 & track_2_3_chanY_n13;
	track_3_2_chanX_n15_driver_mux_fanins <= CLB_3_3_OUT_pin_0 & track_3_2_chanY_n12 & track_4_2_chanX_n15 & track_3_3_chanY_n3;
	track_3_2_chanX_n2_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_2_2_chanY_n10 & track_2_2_chanX_n2 & track_2_3_chanY_n1;
	track_3_2_chanX_n3_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_3_2_chanY_n0 & track_4_2_chanX_n3 & track_3_3_chanY_n15;
	track_3_2_chanX_n4_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_2_2_chanY_n8 & track_2_2_chanX_n4 & track_2_3_chanY_n3;
	track_3_2_chanX_n5_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_3_2_chanY_n2 & track_4_2_chanX_n5 & track_3_3_chanY_n13;
	track_3_2_chanX_n6_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_2_2_chanY_n6 & track_2_2_chanX_n6 & track_2_3_chanY_n5;
	track_3_2_chanX_n7_driver_mux_fanins  <= CLB_3_2_OUT_pin_2 & track_3_2_chanY_n4 & track_4_2_chanX_n7 & track_3_3_chanY_n11;
	track_3_2_chanX_n8_driver_mux_fanins  <= CLB_3_3_OUT_pin_0 & track_2_2_chanY_n4 & track_2_2_chanX_n8 & track_2_3_chanY_n7;
	track_3_2_chanX_n9_driver_mux_fanins  <= CLB_3_3_OUT_pin_0 & track_3_2_chanY_n6 & track_4_2_chanX_n9 & track_3_3_chanY_n9;
	track_3_2_chanY_n0_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_3_1_chanY_n0 & track_4_1_chanX_n3 & track_3_1_chanX_n0;
	track_3_2_chanY_n1_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_4_2_chanX_n13 & track_3_2_chanX_n2 & track_3_3_chanY_n1;
	track_3_2_chanY_n10_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_3_1_chanY_n10 & track_4_1_chanX_n13 & track_3_1_chanX_n6;
	track_3_2_chanY_n11_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_4_2_chanX_n3 & track_3_2_chanX_n12 & track_3_3_chanY_n11;
	track_3_2_chanY_n12_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_3_1_chanY_n12 & track_4_1_chanX_n15 & track_3_1_chanX_n4;
	track_3_2_chanY_n13_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_4_2_chanX_n1 & track_3_2_chanX_n14 & track_3_3_chanY_n13;
	track_3_2_chanY_n14_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_3_1_chanY_n14 & track_4_1_chanX_n1 & track_3_1_chanX_n2;
	track_3_2_chanY_n15_driver_mux_fanins <= CLB_4_2_OUT_pin_1 & track_4_2_chanX_n15 & track_3_2_chanX_n0 & track_3_3_chanY_n15;
	track_3_2_chanY_n2_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_3_1_chanY_n2 & track_4_1_chanX_n5 & track_3_1_chanX_n14;
	track_3_2_chanY_n3_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_4_2_chanX_n11 & track_3_2_chanX_n4 & track_3_3_chanY_n3;
	track_3_2_chanY_n4_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_3_1_chanY_n4 & track_4_1_chanX_n7 & track_3_1_chanX_n12;
	track_3_2_chanY_n5_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_4_2_chanX_n9 & track_3_2_chanX_n6 & track_3_3_chanY_n5;
	track_3_2_chanY_n6_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_3_1_chanY_n6 & track_4_1_chanX_n9 & track_3_1_chanX_n10;
	track_3_2_chanY_n7_driver_mux_fanins  <= CLB_3_2_OUT_pin_3 & track_4_2_chanX_n7 & track_3_2_chanX_n8 & track_3_3_chanY_n7;
	track_3_2_chanY_n8_driver_mux_fanins  <= CLB_4_2_OUT_pin_1 & track_3_1_chanY_n8 & track_4_1_chanX_n11 & track_3_1_chanX_n8;
	track_3_2_chanY_n9_driver_mux_fanins  <= CLB_4_2_OUT_pin_1 & track_4_2_chanX_n5 & track_3_2_chanX_n10 & track_3_3_chanY_n9;
	track_3_3_chanX_n0_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_2_3_chanY_n12 & track_2_3_chanX_n0 & track_2_4_chanY_n15;
	track_3_3_chanX_n1_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_3_3_chanY_n14 & track_4_3_chanX_n1 & track_3_4_chanY_n1;
	track_3_3_chanX_n10_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_2_3_chanY_n2 & track_2_3_chanX_n10 & track_2_4_chanY_n9;
	track_3_3_chanX_n11_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_3_3_chanY_n8 & track_4_3_chanX_n11 & track_3_4_chanY_n7;
	track_3_3_chanX_n12_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_2_3_chanY_n0 & track_2_3_chanX_n12 & track_2_4_chanY_n11;
	track_3_3_chanX_n13_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_3_3_chanY_n10 & track_4_3_chanX_n13 & track_3_4_chanY_n5;
	track_3_3_chanX_n14_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_2_3_chanY_n14 & track_2_3_chanX_n14 & track_2_4_chanY_n13;
	track_3_3_chanX_n15_driver_mux_fanins <= CLB_3_4_OUT_pin_0 & track_3_3_chanY_n12 & track_4_3_chanX_n15 & track_3_4_chanY_n3;
	track_3_3_chanX_n2_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_2_3_chanY_n10 & track_2_3_chanX_n2 & track_2_4_chanY_n1;
	track_3_3_chanX_n3_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_3_3_chanY_n0 & track_4_3_chanX_n3 & track_3_4_chanY_n15;
	track_3_3_chanX_n4_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_2_3_chanY_n8 & track_2_3_chanX_n4 & track_2_4_chanY_n3;
	track_3_3_chanX_n5_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_3_3_chanY_n2 & track_4_3_chanX_n5 & track_3_4_chanY_n13;
	track_3_3_chanX_n6_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_2_3_chanY_n6 & track_2_3_chanX_n6 & track_2_4_chanY_n5;
	track_3_3_chanX_n7_driver_mux_fanins  <= CLB_3_3_OUT_pin_2 & track_3_3_chanY_n4 & track_4_3_chanX_n7 & track_3_4_chanY_n11;
	track_3_3_chanX_n8_driver_mux_fanins  <= CLB_3_4_OUT_pin_0 & track_2_3_chanY_n4 & track_2_3_chanX_n8 & track_2_4_chanY_n7;
	track_3_3_chanX_n9_driver_mux_fanins  <= CLB_3_4_OUT_pin_0 & track_3_3_chanY_n6 & track_4_3_chanX_n9 & track_3_4_chanY_n9;
	track_3_3_chanY_n0_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_3_2_chanY_n0 & track_4_2_chanX_n3 & track_3_2_chanX_n0;
	track_3_3_chanY_n1_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_4_3_chanX_n13 & track_3_3_chanX_n2 & track_3_4_chanY_n1;
	track_3_3_chanY_n10_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_3_2_chanY_n10 & track_4_2_chanX_n13 & track_3_2_chanX_n6;
	track_3_3_chanY_n11_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_4_3_chanX_n3 & track_3_3_chanX_n12 & track_3_4_chanY_n11;
	track_3_3_chanY_n12_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_3_2_chanY_n12 & track_4_2_chanX_n15 & track_3_2_chanX_n4;
	track_3_3_chanY_n13_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_4_3_chanX_n1 & track_3_3_chanX_n14 & track_3_4_chanY_n13;
	track_3_3_chanY_n14_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_3_2_chanY_n14 & track_4_2_chanX_n1 & track_3_2_chanX_n2;
	track_3_3_chanY_n15_driver_mux_fanins <= CLB_4_3_OUT_pin_1 & track_4_3_chanX_n15 & track_3_3_chanX_n0 & track_3_4_chanY_n15;
	track_3_3_chanY_n2_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_3_2_chanY_n2 & track_4_2_chanX_n5 & track_3_2_chanX_n14;
	track_3_3_chanY_n3_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_4_3_chanX_n11 & track_3_3_chanX_n4 & track_3_4_chanY_n3;
	track_3_3_chanY_n4_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_3_2_chanY_n4 & track_4_2_chanX_n7 & track_3_2_chanX_n12;
	track_3_3_chanY_n5_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_4_3_chanX_n9 & track_3_3_chanX_n6 & track_3_4_chanY_n5;
	track_3_3_chanY_n6_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_3_2_chanY_n6 & track_4_2_chanX_n9 & track_3_2_chanX_n10;
	track_3_3_chanY_n7_driver_mux_fanins  <= CLB_3_3_OUT_pin_3 & track_4_3_chanX_n7 & track_3_3_chanX_n8 & track_3_4_chanY_n7;
	track_3_3_chanY_n8_driver_mux_fanins  <= CLB_4_3_OUT_pin_1 & track_3_2_chanY_n8 & track_4_2_chanX_n11 & track_3_2_chanX_n8;
	track_3_3_chanY_n9_driver_mux_fanins  <= CLB_4_3_OUT_pin_1 & track_4_3_chanX_n5 & track_3_3_chanX_n10 & track_3_4_chanY_n9;
	track_3_4_chanX_n0_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_2_4_chanY_n12 & track_2_4_chanX_n0 & track_2_5_chanY_n15;
	track_3_4_chanX_n1_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_3_4_chanY_n14 & track_4_4_chanX_n1 & track_3_5_chanY_n1;
	track_3_4_chanX_n10_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_2_4_chanY_n2 & track_2_4_chanX_n10 & track_2_5_chanY_n9;
	track_3_4_chanX_n11_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_3_4_chanY_n8 & track_4_4_chanX_n11 & track_3_5_chanY_n7;
	track_3_4_chanX_n12_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_2_4_chanY_n0 & track_2_4_chanX_n12 & track_2_5_chanY_n11;
	track_3_4_chanX_n13_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_3_4_chanY_n10 & track_4_4_chanX_n13 & track_3_5_chanY_n5;
	track_3_4_chanX_n14_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_2_4_chanY_n14 & track_2_4_chanX_n14 & track_2_5_chanY_n13;
	track_3_4_chanX_n15_driver_mux_fanins <= CLB_3_5_OUT_pin_0 & track_3_4_chanY_n12 & track_4_4_chanX_n15 & track_3_5_chanY_n3;
	track_3_4_chanX_n2_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_2_4_chanY_n10 & track_2_4_chanX_n2 & track_2_5_chanY_n1;
	track_3_4_chanX_n3_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_3_4_chanY_n0 & track_4_4_chanX_n3 & track_3_5_chanY_n15;
	track_3_4_chanX_n4_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_2_4_chanY_n8 & track_2_4_chanX_n4 & track_2_5_chanY_n3;
	track_3_4_chanX_n5_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_3_4_chanY_n2 & track_4_4_chanX_n5 & track_3_5_chanY_n13;
	track_3_4_chanX_n6_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_2_4_chanY_n6 & track_2_4_chanX_n6 & track_2_5_chanY_n5;
	track_3_4_chanX_n7_driver_mux_fanins  <= CLB_3_4_OUT_pin_2 & track_3_4_chanY_n4 & track_4_4_chanX_n7 & track_3_5_chanY_n11;
	track_3_4_chanX_n8_driver_mux_fanins  <= CLB_3_5_OUT_pin_0 & track_2_4_chanY_n4 & track_2_4_chanX_n8 & track_2_5_chanY_n7;
	track_3_4_chanX_n9_driver_mux_fanins  <= CLB_3_5_OUT_pin_0 & track_3_4_chanY_n6 & track_4_4_chanX_n9 & track_3_5_chanY_n9;
	track_3_4_chanY_n0_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_3_3_chanY_n0 & track_4_3_chanX_n3 & track_3_3_chanX_n0;
	track_3_4_chanY_n1_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_4_4_chanX_n13 & track_3_4_chanX_n2 & track_3_5_chanY_n1;
	track_3_4_chanY_n10_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_3_3_chanY_n10 & track_4_3_chanX_n13 & track_3_3_chanX_n6;
	track_3_4_chanY_n11_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_4_4_chanX_n3 & track_3_4_chanX_n12 & track_3_5_chanY_n11;
	track_3_4_chanY_n12_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_3_3_chanY_n12 & track_4_3_chanX_n15 & track_3_3_chanX_n4;
	track_3_4_chanY_n13_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_4_4_chanX_n1 & track_3_4_chanX_n14 & track_3_5_chanY_n13;
	track_3_4_chanY_n14_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_3_3_chanY_n14 & track_4_3_chanX_n1 & track_3_3_chanX_n2;
	track_3_4_chanY_n15_driver_mux_fanins <= CLB_4_4_OUT_pin_1 & track_4_4_chanX_n15 & track_3_4_chanX_n0 & track_3_5_chanY_n15;
	track_3_4_chanY_n2_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_3_3_chanY_n2 & track_4_3_chanX_n5 & track_3_3_chanX_n14;
	track_3_4_chanY_n3_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_4_4_chanX_n11 & track_3_4_chanX_n4 & track_3_5_chanY_n3;
	track_3_4_chanY_n4_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_3_3_chanY_n4 & track_4_3_chanX_n7 & track_3_3_chanX_n12;
	track_3_4_chanY_n5_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_4_4_chanX_n9 & track_3_4_chanX_n6 & track_3_5_chanY_n5;
	track_3_4_chanY_n6_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_3_3_chanY_n6 & track_4_3_chanX_n9 & track_3_3_chanX_n10;
	track_3_4_chanY_n7_driver_mux_fanins  <= CLB_3_4_OUT_pin_3 & track_4_4_chanX_n7 & track_3_4_chanX_n8 & track_3_5_chanY_n7;
	track_3_4_chanY_n8_driver_mux_fanins  <= CLB_4_4_OUT_pin_1 & track_3_3_chanY_n8 & track_4_3_chanX_n11 & track_3_3_chanX_n8;
	track_3_4_chanY_n9_driver_mux_fanins  <= CLB_4_4_OUT_pin_1 & track_4_4_chanX_n5 & track_3_4_chanX_n10 & track_3_5_chanY_n9;
	track_3_5_chanX_n0_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_2_5_chanY_n12 & track_2_5_chanX_n0 & track_2_6_chanY_n15;
	track_3_5_chanX_n1_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_3_5_chanY_n14 & track_4_5_chanX_n1 & track_3_6_chanY_n1;
	track_3_5_chanX_n10_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_2_5_chanY_n2 & track_2_5_chanX_n10 & track_2_6_chanY_n9;
	track_3_5_chanX_n11_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_3_5_chanY_n8 & track_4_5_chanX_n11 & track_3_6_chanY_n7;
	track_3_5_chanX_n12_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_2_5_chanY_n0 & track_2_5_chanX_n12 & track_2_6_chanY_n11;
	track_3_5_chanX_n13_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_3_5_chanY_n10 & track_4_5_chanX_n13 & track_3_6_chanY_n5;
	track_3_5_chanX_n14_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_2_5_chanY_n14 & track_2_5_chanX_n14 & track_2_6_chanY_n13;
	track_3_5_chanX_n15_driver_mux_fanins <= CLB_3_6_OUT_pin_0 & track_3_5_chanY_n12 & track_4_5_chanX_n15 & track_3_6_chanY_n3;
	track_3_5_chanX_n2_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_2_5_chanY_n10 & track_2_5_chanX_n2 & track_2_6_chanY_n1;
	track_3_5_chanX_n3_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_3_5_chanY_n0 & track_4_5_chanX_n3 & track_3_6_chanY_n15;
	track_3_5_chanX_n4_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_2_5_chanY_n8 & track_2_5_chanX_n4 & track_2_6_chanY_n3;
	track_3_5_chanX_n5_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_3_5_chanY_n2 & track_4_5_chanX_n5 & track_3_6_chanY_n13;
	track_3_5_chanX_n6_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_2_5_chanY_n6 & track_2_5_chanX_n6 & track_2_6_chanY_n5;
	track_3_5_chanX_n7_driver_mux_fanins  <= CLB_3_5_OUT_pin_2 & track_3_5_chanY_n4 & track_4_5_chanX_n7 & track_3_6_chanY_n11;
	track_3_5_chanX_n8_driver_mux_fanins  <= CLB_3_6_OUT_pin_0 & track_2_5_chanY_n4 & track_2_5_chanX_n8 & track_2_6_chanY_n7;
	track_3_5_chanX_n9_driver_mux_fanins  <= CLB_3_6_OUT_pin_0 & track_3_5_chanY_n6 & track_4_5_chanX_n9 & track_3_6_chanY_n9;
	track_3_5_chanY_n0_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_3_4_chanY_n0 & track_4_4_chanX_n3 & track_3_4_chanX_n0;
	track_3_5_chanY_n1_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_4_5_chanX_n13 & track_3_5_chanX_n2 & track_3_6_chanY_n1;
	track_3_5_chanY_n10_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_3_4_chanY_n10 & track_4_4_chanX_n13 & track_3_4_chanX_n6;
	track_3_5_chanY_n11_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_4_5_chanX_n3 & track_3_5_chanX_n12 & track_3_6_chanY_n11;
	track_3_5_chanY_n12_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_3_4_chanY_n12 & track_4_4_chanX_n15 & track_3_4_chanX_n4;
	track_3_5_chanY_n13_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_4_5_chanX_n1 & track_3_5_chanX_n14 & track_3_6_chanY_n13;
	track_3_5_chanY_n14_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_3_4_chanY_n14 & track_4_4_chanX_n1 & track_3_4_chanX_n2;
	track_3_5_chanY_n15_driver_mux_fanins <= CLB_4_5_OUT_pin_1 & track_4_5_chanX_n15 & track_3_5_chanX_n0 & track_3_6_chanY_n15;
	track_3_5_chanY_n2_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_3_4_chanY_n2 & track_4_4_chanX_n5 & track_3_4_chanX_n14;
	track_3_5_chanY_n3_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_4_5_chanX_n11 & track_3_5_chanX_n4 & track_3_6_chanY_n3;
	track_3_5_chanY_n4_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_3_4_chanY_n4 & track_4_4_chanX_n7 & track_3_4_chanX_n12;
	track_3_5_chanY_n5_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_4_5_chanX_n9 & track_3_5_chanX_n6 & track_3_6_chanY_n5;
	track_3_5_chanY_n6_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_3_4_chanY_n6 & track_4_4_chanX_n9 & track_3_4_chanX_n10;
	track_3_5_chanY_n7_driver_mux_fanins  <= CLB_3_5_OUT_pin_3 & track_4_5_chanX_n7 & track_3_5_chanX_n8 & track_3_6_chanY_n7;
	track_3_5_chanY_n8_driver_mux_fanins  <= CLB_4_5_OUT_pin_1 & track_3_4_chanY_n8 & track_4_4_chanX_n11 & track_3_4_chanX_n8;
	track_3_5_chanY_n9_driver_mux_fanins  <= CLB_4_5_OUT_pin_1 & track_4_5_chanX_n5 & track_3_5_chanX_n10 & track_3_6_chanY_n9;
	track_3_6_chanX_n0_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_2_6_chanY_n0 & track_2_6_chanX_n0;
	track_3_6_chanX_n1_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_3_6_chanY_n0 & track_4_6_chanX_n1;
	track_3_6_chanX_n10_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_2_6_chanY_n10 & track_2_6_chanX_n10;
	track_3_6_chanX_n11_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_3_6_chanY_n10 & track_4_6_chanX_n11;
	track_3_6_chanX_n12_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_2_6_chanY_n12 & track_2_6_chanX_n12;
	track_3_6_chanX_n13_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_3_6_chanY_n12 & track_4_6_chanX_n13;
	track_3_6_chanX_n14_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_2_6_chanY_n14 & track_2_6_chanX_n14;
	track_3_6_chanX_n15_driver_mux_fanins <= "0" & IO_3_7_OUT_pin_0 & track_3_6_chanY_n14 & track_4_6_chanX_n15;
	track_3_6_chanX_n2_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_2_6_chanY_n2 & track_2_6_chanX_n2;
	track_3_6_chanX_n3_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_3_6_chanY_n2 & track_4_6_chanX_n3;
	track_3_6_chanX_n4_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_2_6_chanY_n4 & track_2_6_chanX_n4;
	track_3_6_chanX_n5_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_3_6_chanY_n4 & track_4_6_chanX_n5;
	track_3_6_chanX_n6_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_2_6_chanY_n6 & track_2_6_chanX_n6;
	track_3_6_chanX_n7_driver_mux_fanins  <= IO_3_7_OUT_pin_1 & CLB_3_6_OUT_pin_2 & track_3_6_chanY_n6 & track_4_6_chanX_n7;
	track_3_6_chanX_n8_driver_mux_fanins  <= "0" & IO_3_7_OUT_pin_0 & track_2_6_chanY_n8 & track_2_6_chanX_n8;
	track_3_6_chanX_n9_driver_mux_fanins  <= "0" & IO_3_7_OUT_pin_0 & track_3_6_chanY_n8 & track_4_6_chanX_n9;
	track_3_6_chanY_n0_driver_mux_fanins  <= CLB_3_6_OUT_pin_3 & track_3_5_chanY_n0 & track_4_5_chanX_n3 & track_3_5_chanX_n0;
	track_3_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_3_6_OUT_pin_3 & track_4_6_chanX_n1 & track_3_6_chanX_n0;
	track_3_6_chanY_n10_driver_mux_fanins <= CLB_4_6_OUT_pin_1 & track_3_5_chanY_n10 & track_4_5_chanX_n13 & track_3_5_chanX_n6;
	track_3_6_chanY_n11_driver_mux_fanins <= "0" & CLB_4_6_OUT_pin_1 & track_4_6_chanX_n5 & track_3_6_chanX_n4;
	track_3_6_chanY_n12_driver_mux_fanins <= CLB_4_6_OUT_pin_1 & track_3_5_chanY_n12 & track_4_5_chanX_n15 & track_3_5_chanX_n4;
	track_3_6_chanY_n13_driver_mux_fanins <= "0" & CLB_4_6_OUT_pin_1 & track_4_6_chanX_n7 & track_3_6_chanX_n6;
	track_3_6_chanY_n14_driver_mux_fanins <= CLB_4_6_OUT_pin_1 & track_3_5_chanY_n14 & track_4_5_chanX_n1 & track_3_5_chanX_n2;
	track_3_6_chanY_n15_driver_mux_fanins <= "0" & CLB_4_6_OUT_pin_1 & track_4_6_chanX_n15 & track_3_6_chanX_n14;
	track_3_6_chanY_n2_driver_mux_fanins  <= CLB_3_6_OUT_pin_3 & track_3_5_chanY_n2 & track_4_5_chanX_n5 & track_3_5_chanX_n14;
	track_3_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_3_6_OUT_pin_3 & track_4_6_chanX_n9 & track_3_6_chanX_n8;
	track_3_6_chanY_n4_driver_mux_fanins  <= CLB_3_6_OUT_pin_3 & track_3_5_chanY_n4 & track_4_5_chanX_n7 & track_3_5_chanX_n12;
	track_3_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_3_6_OUT_pin_3 & track_4_6_chanX_n11 & track_3_6_chanX_n10;
	track_3_6_chanY_n6_driver_mux_fanins  <= CLB_3_6_OUT_pin_3 & track_3_5_chanY_n6 & track_4_5_chanX_n9 & track_3_5_chanX_n10;
	track_3_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_3_6_OUT_pin_3 & track_4_6_chanX_n13 & track_3_6_chanX_n12;
	track_3_6_chanY_n8_driver_mux_fanins  <= CLB_4_6_OUT_pin_1 & track_3_5_chanY_n8 & track_4_5_chanX_n11 & track_3_5_chanX_n8;
	track_3_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_4_6_OUT_pin_1 & track_4_6_chanX_n3 & track_3_6_chanX_n2;
	track_4_0_chanX_n0_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_3_0_chanX_n0 & track_3_1_chanY_n1;
	track_4_0_chanX_n1_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_5_0_chanX_n1 & track_4_1_chanY_n1;
	track_4_0_chanX_n10_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_3_0_chanX_n10 & track_3_1_chanY_n11;
	track_4_0_chanX_n11_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_5_0_chanX_n11 & track_4_1_chanY_n11;
	track_4_0_chanX_n12_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_3_0_chanX_n12 & track_3_1_chanY_n13;
	track_4_0_chanX_n13_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_5_0_chanX_n13 & track_4_1_chanY_n13;
	track_4_0_chanX_n14_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_3_0_chanX_n14 & track_3_1_chanY_n15;
	track_4_0_chanX_n15_driver_mux_fanins <= "0" & IO_4_0_OUT_pin_1 & track_5_0_chanX_n15 & track_4_1_chanY_n15;
	track_4_0_chanX_n2_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_3_0_chanX_n2 & track_3_1_chanY_n3;
	track_4_0_chanX_n3_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_5_0_chanX_n3 & track_4_1_chanY_n3;
	track_4_0_chanX_n4_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_3_0_chanX_n4 & track_3_1_chanY_n5;
	track_4_0_chanX_n5_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_5_0_chanX_n5 & track_4_1_chanY_n5;
	track_4_0_chanX_n6_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_3_0_chanX_n6 & track_3_1_chanY_n7;
	track_4_0_chanX_n7_driver_mux_fanins  <= IO_4_0_OUT_pin_0 & CLB_4_1_OUT_pin_0 & track_5_0_chanX_n7 & track_4_1_chanY_n7;
	track_4_0_chanX_n8_driver_mux_fanins  <= "0" & IO_4_0_OUT_pin_1 & track_3_0_chanX_n8 & track_3_1_chanY_n9;
	track_4_0_chanX_n9_driver_mux_fanins  <= "0" & IO_4_0_OUT_pin_1 & track_5_0_chanX_n9 & track_4_1_chanY_n9;
	track_4_1_chanX_n0_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_3_1_chanY_n12 & track_3_1_chanX_n0 & track_3_2_chanY_n15;
	track_4_1_chanX_n1_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_4_1_chanY_n14 & track_5_1_chanX_n1 & track_4_2_chanY_n1;
	track_4_1_chanX_n10_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_3_1_chanY_n2 & track_3_1_chanX_n10 & track_3_2_chanY_n9;
	track_4_1_chanX_n11_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_4_1_chanY_n8 & track_5_1_chanX_n11 & track_4_2_chanY_n7;
	track_4_1_chanX_n12_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_3_1_chanY_n0 & track_3_1_chanX_n12 & track_3_2_chanY_n11;
	track_4_1_chanX_n13_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_4_1_chanY_n10 & track_5_1_chanX_n13 & track_4_2_chanY_n5;
	track_4_1_chanX_n14_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_3_1_chanY_n14 & track_3_1_chanX_n14 & track_3_2_chanY_n13;
	track_4_1_chanX_n15_driver_mux_fanins <= CLB_4_2_OUT_pin_0 & track_4_1_chanY_n12 & track_5_1_chanX_n15 & track_4_2_chanY_n3;
	track_4_1_chanX_n2_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_3_1_chanY_n10 & track_3_1_chanX_n2 & track_3_2_chanY_n1;
	track_4_1_chanX_n3_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_4_1_chanY_n0 & track_5_1_chanX_n3 & track_4_2_chanY_n15;
	track_4_1_chanX_n4_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_3_1_chanY_n8 & track_3_1_chanX_n4 & track_3_2_chanY_n3;
	track_4_1_chanX_n5_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_4_1_chanY_n2 & track_5_1_chanX_n5 & track_4_2_chanY_n13;
	track_4_1_chanX_n6_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_3_1_chanY_n6 & track_3_1_chanX_n6 & track_3_2_chanY_n5;
	track_4_1_chanX_n7_driver_mux_fanins  <= CLB_4_1_OUT_pin_2 & track_4_1_chanY_n4 & track_5_1_chanX_n7 & track_4_2_chanY_n11;
	track_4_1_chanX_n8_driver_mux_fanins  <= CLB_4_2_OUT_pin_0 & track_3_1_chanY_n4 & track_3_1_chanX_n8 & track_3_2_chanY_n7;
	track_4_1_chanX_n9_driver_mux_fanins  <= CLB_4_2_OUT_pin_0 & track_4_1_chanY_n6 & track_5_1_chanX_n9 & track_4_2_chanY_n9;
	track_4_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_4_1_OUT_pin_3 & track_5_0_chanX_n7 & track_4_0_chanX_n6;
	track_4_1_chanY_n1_driver_mux_fanins  <= CLB_4_1_OUT_pin_3 & track_5_1_chanX_n13 & track_4_1_chanX_n2 & track_4_2_chanY_n1;
	track_4_1_chanY_n10_driver_mux_fanins <= "0" & CLB_5_1_OUT_pin_1 & track_5_0_chanX_n11 & track_4_0_chanX_n10;
	track_4_1_chanY_n11_driver_mux_fanins <= CLB_5_1_OUT_pin_1 & track_5_1_chanX_n3 & track_4_1_chanX_n12 & track_4_2_chanY_n11;
	track_4_1_chanY_n12_driver_mux_fanins <= "0" & CLB_5_1_OUT_pin_1 & track_5_0_chanX_n13 & track_4_0_chanX_n12;
	track_4_1_chanY_n13_driver_mux_fanins <= CLB_5_1_OUT_pin_1 & track_5_1_chanX_n1 & track_4_1_chanX_n14 & track_4_2_chanY_n13;
	track_4_1_chanY_n14_driver_mux_fanins <= "0" & CLB_5_1_OUT_pin_1 & track_5_0_chanX_n15 & track_4_0_chanX_n14;
	track_4_1_chanY_n15_driver_mux_fanins <= CLB_5_1_OUT_pin_1 & track_5_1_chanX_n15 & track_4_1_chanX_n0 & track_4_2_chanY_n15;
	track_4_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_4_1_OUT_pin_3 & track_5_0_chanX_n9 & track_4_0_chanX_n8;
	track_4_1_chanY_n3_driver_mux_fanins  <= CLB_4_1_OUT_pin_3 & track_5_1_chanX_n11 & track_4_1_chanX_n4 & track_4_2_chanY_n3;
	track_4_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_4_1_OUT_pin_3 & track_5_0_chanX_n1 & track_4_0_chanX_n0;
	track_4_1_chanY_n5_driver_mux_fanins  <= CLB_4_1_OUT_pin_3 & track_5_1_chanX_n9 & track_4_1_chanX_n6 & track_4_2_chanY_n5;
	track_4_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_4_1_OUT_pin_3 & track_5_0_chanX_n3 & track_4_0_chanX_n2;
	track_4_1_chanY_n7_driver_mux_fanins  <= CLB_4_1_OUT_pin_3 & track_5_1_chanX_n7 & track_4_1_chanX_n8 & track_4_2_chanY_n7;
	track_4_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_5_1_OUT_pin_1 & track_5_0_chanX_n5 & track_4_0_chanX_n4;
	track_4_1_chanY_n9_driver_mux_fanins  <= CLB_5_1_OUT_pin_1 & track_5_1_chanX_n5 & track_4_1_chanX_n10 & track_4_2_chanY_n9;
	track_4_2_chanX_n0_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_3_2_chanY_n12 & track_3_2_chanX_n0 & track_3_3_chanY_n15;
	track_4_2_chanX_n1_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_4_2_chanY_n14 & track_5_2_chanX_n1 & track_4_3_chanY_n1;
	track_4_2_chanX_n10_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_3_2_chanY_n2 & track_3_2_chanX_n10 & track_3_3_chanY_n9;
	track_4_2_chanX_n11_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_4_2_chanY_n8 & track_5_2_chanX_n11 & track_4_3_chanY_n7;
	track_4_2_chanX_n12_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_3_2_chanY_n0 & track_3_2_chanX_n12 & track_3_3_chanY_n11;
	track_4_2_chanX_n13_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_4_2_chanY_n10 & track_5_2_chanX_n13 & track_4_3_chanY_n5;
	track_4_2_chanX_n14_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_3_2_chanY_n14 & track_3_2_chanX_n14 & track_3_3_chanY_n13;
	track_4_2_chanX_n15_driver_mux_fanins <= CLB_4_3_OUT_pin_0 & track_4_2_chanY_n12 & track_5_2_chanX_n15 & track_4_3_chanY_n3;
	track_4_2_chanX_n2_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_3_2_chanY_n10 & track_3_2_chanX_n2 & track_3_3_chanY_n1;
	track_4_2_chanX_n3_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_4_2_chanY_n0 & track_5_2_chanX_n3 & track_4_3_chanY_n15;
	track_4_2_chanX_n4_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_3_2_chanY_n8 & track_3_2_chanX_n4 & track_3_3_chanY_n3;
	track_4_2_chanX_n5_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_4_2_chanY_n2 & track_5_2_chanX_n5 & track_4_3_chanY_n13;
	track_4_2_chanX_n6_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_3_2_chanY_n6 & track_3_2_chanX_n6 & track_3_3_chanY_n5;
	track_4_2_chanX_n7_driver_mux_fanins  <= CLB_4_2_OUT_pin_2 & track_4_2_chanY_n4 & track_5_2_chanX_n7 & track_4_3_chanY_n11;
	track_4_2_chanX_n8_driver_mux_fanins  <= CLB_4_3_OUT_pin_0 & track_3_2_chanY_n4 & track_3_2_chanX_n8 & track_3_3_chanY_n7;
	track_4_2_chanX_n9_driver_mux_fanins  <= CLB_4_3_OUT_pin_0 & track_4_2_chanY_n6 & track_5_2_chanX_n9 & track_4_3_chanY_n9;
	track_4_2_chanY_n0_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_4_1_chanY_n0 & track_5_1_chanX_n3 & track_4_1_chanX_n0;
	track_4_2_chanY_n1_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_5_2_chanX_n13 & track_4_2_chanX_n2 & track_4_3_chanY_n1;
	track_4_2_chanY_n10_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_4_1_chanY_n10 & track_5_1_chanX_n13 & track_4_1_chanX_n6;
	track_4_2_chanY_n11_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_5_2_chanX_n3 & track_4_2_chanX_n12 & track_4_3_chanY_n11;
	track_4_2_chanY_n12_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_4_1_chanY_n12 & track_5_1_chanX_n15 & track_4_1_chanX_n4;
	track_4_2_chanY_n13_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_5_2_chanX_n1 & track_4_2_chanX_n14 & track_4_3_chanY_n13;
	track_4_2_chanY_n14_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_4_1_chanY_n14 & track_5_1_chanX_n1 & track_4_1_chanX_n2;
	track_4_2_chanY_n15_driver_mux_fanins <= CLB_5_2_OUT_pin_1 & track_5_2_chanX_n15 & track_4_2_chanX_n0 & track_4_3_chanY_n15;
	track_4_2_chanY_n2_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_4_1_chanY_n2 & track_5_1_chanX_n5 & track_4_1_chanX_n14;
	track_4_2_chanY_n3_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_5_2_chanX_n11 & track_4_2_chanX_n4 & track_4_3_chanY_n3;
	track_4_2_chanY_n4_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_4_1_chanY_n4 & track_5_1_chanX_n7 & track_4_1_chanX_n12;
	track_4_2_chanY_n5_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_5_2_chanX_n9 & track_4_2_chanX_n6 & track_4_3_chanY_n5;
	track_4_2_chanY_n6_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_4_1_chanY_n6 & track_5_1_chanX_n9 & track_4_1_chanX_n10;
	track_4_2_chanY_n7_driver_mux_fanins  <= CLB_4_2_OUT_pin_3 & track_5_2_chanX_n7 & track_4_2_chanX_n8 & track_4_3_chanY_n7;
	track_4_2_chanY_n8_driver_mux_fanins  <= CLB_5_2_OUT_pin_1 & track_4_1_chanY_n8 & track_5_1_chanX_n11 & track_4_1_chanX_n8;
	track_4_2_chanY_n9_driver_mux_fanins  <= CLB_5_2_OUT_pin_1 & track_5_2_chanX_n5 & track_4_2_chanX_n10 & track_4_3_chanY_n9;
	track_4_3_chanX_n0_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_3_3_chanY_n12 & track_3_3_chanX_n0 & track_3_4_chanY_n15;
	track_4_3_chanX_n1_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_4_3_chanY_n14 & track_5_3_chanX_n1 & track_4_4_chanY_n1;
	track_4_3_chanX_n10_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_3_3_chanY_n2 & track_3_3_chanX_n10 & track_3_4_chanY_n9;
	track_4_3_chanX_n11_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_4_3_chanY_n8 & track_5_3_chanX_n11 & track_4_4_chanY_n7;
	track_4_3_chanX_n12_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_3_3_chanY_n0 & track_3_3_chanX_n12 & track_3_4_chanY_n11;
	track_4_3_chanX_n13_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_4_3_chanY_n10 & track_5_3_chanX_n13 & track_4_4_chanY_n5;
	track_4_3_chanX_n14_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_3_3_chanY_n14 & track_3_3_chanX_n14 & track_3_4_chanY_n13;
	track_4_3_chanX_n15_driver_mux_fanins <= CLB_4_4_OUT_pin_0 & track_4_3_chanY_n12 & track_5_3_chanX_n15 & track_4_4_chanY_n3;
	track_4_3_chanX_n2_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_3_3_chanY_n10 & track_3_3_chanX_n2 & track_3_4_chanY_n1;
	track_4_3_chanX_n3_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_4_3_chanY_n0 & track_5_3_chanX_n3 & track_4_4_chanY_n15;
	track_4_3_chanX_n4_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_3_3_chanY_n8 & track_3_3_chanX_n4 & track_3_4_chanY_n3;
	track_4_3_chanX_n5_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_4_3_chanY_n2 & track_5_3_chanX_n5 & track_4_4_chanY_n13;
	track_4_3_chanX_n6_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_3_3_chanY_n6 & track_3_3_chanX_n6 & track_3_4_chanY_n5;
	track_4_3_chanX_n7_driver_mux_fanins  <= CLB_4_3_OUT_pin_2 & track_4_3_chanY_n4 & track_5_3_chanX_n7 & track_4_4_chanY_n11;
	track_4_3_chanX_n8_driver_mux_fanins  <= CLB_4_4_OUT_pin_0 & track_3_3_chanY_n4 & track_3_3_chanX_n8 & track_3_4_chanY_n7;
	track_4_3_chanX_n9_driver_mux_fanins  <= CLB_4_4_OUT_pin_0 & track_4_3_chanY_n6 & track_5_3_chanX_n9 & track_4_4_chanY_n9;
	track_4_3_chanY_n0_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_4_2_chanY_n0 & track_5_2_chanX_n3 & track_4_2_chanX_n0;
	track_4_3_chanY_n1_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_5_3_chanX_n13 & track_4_3_chanX_n2 & track_4_4_chanY_n1;
	track_4_3_chanY_n10_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_4_2_chanY_n10 & track_5_2_chanX_n13 & track_4_2_chanX_n6;
	track_4_3_chanY_n11_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_5_3_chanX_n3 & track_4_3_chanX_n12 & track_4_4_chanY_n11;
	track_4_3_chanY_n12_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_4_2_chanY_n12 & track_5_2_chanX_n15 & track_4_2_chanX_n4;
	track_4_3_chanY_n13_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_5_3_chanX_n1 & track_4_3_chanX_n14 & track_4_4_chanY_n13;
	track_4_3_chanY_n14_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_4_2_chanY_n14 & track_5_2_chanX_n1 & track_4_2_chanX_n2;
	track_4_3_chanY_n15_driver_mux_fanins <= CLB_5_3_OUT_pin_1 & track_5_3_chanX_n15 & track_4_3_chanX_n0 & track_4_4_chanY_n15;
	track_4_3_chanY_n2_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_4_2_chanY_n2 & track_5_2_chanX_n5 & track_4_2_chanX_n14;
	track_4_3_chanY_n3_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_5_3_chanX_n11 & track_4_3_chanX_n4 & track_4_4_chanY_n3;
	track_4_3_chanY_n4_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_4_2_chanY_n4 & track_5_2_chanX_n7 & track_4_2_chanX_n12;
	track_4_3_chanY_n5_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_5_3_chanX_n9 & track_4_3_chanX_n6 & track_4_4_chanY_n5;
	track_4_3_chanY_n6_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_4_2_chanY_n6 & track_5_2_chanX_n9 & track_4_2_chanX_n10;
	track_4_3_chanY_n7_driver_mux_fanins  <= CLB_4_3_OUT_pin_3 & track_5_3_chanX_n7 & track_4_3_chanX_n8 & track_4_4_chanY_n7;
	track_4_3_chanY_n8_driver_mux_fanins  <= CLB_5_3_OUT_pin_1 & track_4_2_chanY_n8 & track_5_2_chanX_n11 & track_4_2_chanX_n8;
	track_4_3_chanY_n9_driver_mux_fanins  <= CLB_5_3_OUT_pin_1 & track_5_3_chanX_n5 & track_4_3_chanX_n10 & track_4_4_chanY_n9;
	track_4_4_chanX_n0_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_3_4_chanY_n12 & track_3_4_chanX_n0 & track_3_5_chanY_n15;
	track_4_4_chanX_n1_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_4_4_chanY_n14 & track_5_4_chanX_n1 & track_4_5_chanY_n1;
	track_4_4_chanX_n10_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_3_4_chanY_n2 & track_3_4_chanX_n10 & track_3_5_chanY_n9;
	track_4_4_chanX_n11_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_4_4_chanY_n8 & track_5_4_chanX_n11 & track_4_5_chanY_n7;
	track_4_4_chanX_n12_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_3_4_chanY_n0 & track_3_4_chanX_n12 & track_3_5_chanY_n11;
	track_4_4_chanX_n13_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_4_4_chanY_n10 & track_5_4_chanX_n13 & track_4_5_chanY_n5;
	track_4_4_chanX_n14_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_3_4_chanY_n14 & track_3_4_chanX_n14 & track_3_5_chanY_n13;
	track_4_4_chanX_n15_driver_mux_fanins <= CLB_4_5_OUT_pin_0 & track_4_4_chanY_n12 & track_5_4_chanX_n15 & track_4_5_chanY_n3;
	track_4_4_chanX_n2_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_3_4_chanY_n10 & track_3_4_chanX_n2 & track_3_5_chanY_n1;
	track_4_4_chanX_n3_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_4_4_chanY_n0 & track_5_4_chanX_n3 & track_4_5_chanY_n15;
	track_4_4_chanX_n4_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_3_4_chanY_n8 & track_3_4_chanX_n4 & track_3_5_chanY_n3;
	track_4_4_chanX_n5_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_4_4_chanY_n2 & track_5_4_chanX_n5 & track_4_5_chanY_n13;
	track_4_4_chanX_n6_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_3_4_chanY_n6 & track_3_4_chanX_n6 & track_3_5_chanY_n5;
	track_4_4_chanX_n7_driver_mux_fanins  <= CLB_4_4_OUT_pin_2 & track_4_4_chanY_n4 & track_5_4_chanX_n7 & track_4_5_chanY_n11;
	track_4_4_chanX_n8_driver_mux_fanins  <= CLB_4_5_OUT_pin_0 & track_3_4_chanY_n4 & track_3_4_chanX_n8 & track_3_5_chanY_n7;
	track_4_4_chanX_n9_driver_mux_fanins  <= CLB_4_5_OUT_pin_0 & track_4_4_chanY_n6 & track_5_4_chanX_n9 & track_4_5_chanY_n9;
	track_4_4_chanY_n0_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_4_3_chanY_n0 & track_5_3_chanX_n3 & track_4_3_chanX_n0;
	track_4_4_chanY_n1_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_5_4_chanX_n13 & track_4_4_chanX_n2 & track_4_5_chanY_n1;
	track_4_4_chanY_n10_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_4_3_chanY_n10 & track_5_3_chanX_n13 & track_4_3_chanX_n6;
	track_4_4_chanY_n11_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_5_4_chanX_n3 & track_4_4_chanX_n12 & track_4_5_chanY_n11;
	track_4_4_chanY_n12_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_4_3_chanY_n12 & track_5_3_chanX_n15 & track_4_3_chanX_n4;
	track_4_4_chanY_n13_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_5_4_chanX_n1 & track_4_4_chanX_n14 & track_4_5_chanY_n13;
	track_4_4_chanY_n14_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_4_3_chanY_n14 & track_5_3_chanX_n1 & track_4_3_chanX_n2;
	track_4_4_chanY_n15_driver_mux_fanins <= CLB_5_4_OUT_pin_1 & track_5_4_chanX_n15 & track_4_4_chanX_n0 & track_4_5_chanY_n15;
	track_4_4_chanY_n2_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_4_3_chanY_n2 & track_5_3_chanX_n5 & track_4_3_chanX_n14;
	track_4_4_chanY_n3_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_5_4_chanX_n11 & track_4_4_chanX_n4 & track_4_5_chanY_n3;
	track_4_4_chanY_n4_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_4_3_chanY_n4 & track_5_3_chanX_n7 & track_4_3_chanX_n12;
	track_4_4_chanY_n5_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_5_4_chanX_n9 & track_4_4_chanX_n6 & track_4_5_chanY_n5;
	track_4_4_chanY_n6_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_4_3_chanY_n6 & track_5_3_chanX_n9 & track_4_3_chanX_n10;
	track_4_4_chanY_n7_driver_mux_fanins  <= CLB_4_4_OUT_pin_3 & track_5_4_chanX_n7 & track_4_4_chanX_n8 & track_4_5_chanY_n7;
	track_4_4_chanY_n8_driver_mux_fanins  <= CLB_5_4_OUT_pin_1 & track_4_3_chanY_n8 & track_5_3_chanX_n11 & track_4_3_chanX_n8;
	track_4_4_chanY_n9_driver_mux_fanins  <= CLB_5_4_OUT_pin_1 & track_5_4_chanX_n5 & track_4_4_chanX_n10 & track_4_5_chanY_n9;
	track_4_5_chanX_n0_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_3_5_chanY_n12 & track_3_5_chanX_n0 & track_3_6_chanY_n15;
	track_4_5_chanX_n1_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_4_5_chanY_n14 & track_5_5_chanX_n1 & track_4_6_chanY_n1;
	track_4_5_chanX_n10_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_3_5_chanY_n2 & track_3_5_chanX_n10 & track_3_6_chanY_n9;
	track_4_5_chanX_n11_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_4_5_chanY_n8 & track_5_5_chanX_n11 & track_4_6_chanY_n7;
	track_4_5_chanX_n12_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_3_5_chanY_n0 & track_3_5_chanX_n12 & track_3_6_chanY_n11;
	track_4_5_chanX_n13_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_4_5_chanY_n10 & track_5_5_chanX_n13 & track_4_6_chanY_n5;
	track_4_5_chanX_n14_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_3_5_chanY_n14 & track_3_5_chanX_n14 & track_3_6_chanY_n13;
	track_4_5_chanX_n15_driver_mux_fanins <= CLB_4_6_OUT_pin_0 & track_4_5_chanY_n12 & track_5_5_chanX_n15 & track_4_6_chanY_n3;
	track_4_5_chanX_n2_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_3_5_chanY_n10 & track_3_5_chanX_n2 & track_3_6_chanY_n1;
	track_4_5_chanX_n3_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_4_5_chanY_n0 & track_5_5_chanX_n3 & track_4_6_chanY_n15;
	track_4_5_chanX_n4_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_3_5_chanY_n8 & track_3_5_chanX_n4 & track_3_6_chanY_n3;
	track_4_5_chanX_n5_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_4_5_chanY_n2 & track_5_5_chanX_n5 & track_4_6_chanY_n13;
	track_4_5_chanX_n6_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_3_5_chanY_n6 & track_3_5_chanX_n6 & track_3_6_chanY_n5;
	track_4_5_chanX_n7_driver_mux_fanins  <= CLB_4_5_OUT_pin_2 & track_4_5_chanY_n4 & track_5_5_chanX_n7 & track_4_6_chanY_n11;
	track_4_5_chanX_n8_driver_mux_fanins  <= CLB_4_6_OUT_pin_0 & track_3_5_chanY_n4 & track_3_5_chanX_n8 & track_3_6_chanY_n7;
	track_4_5_chanX_n9_driver_mux_fanins  <= CLB_4_6_OUT_pin_0 & track_4_5_chanY_n6 & track_5_5_chanX_n9 & track_4_6_chanY_n9;
	track_4_5_chanY_n0_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_4_4_chanY_n0 & track_5_4_chanX_n3 & track_4_4_chanX_n0;
	track_4_5_chanY_n1_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_5_5_chanX_n13 & track_4_5_chanX_n2 & track_4_6_chanY_n1;
	track_4_5_chanY_n10_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_4_4_chanY_n10 & track_5_4_chanX_n13 & track_4_4_chanX_n6;
	track_4_5_chanY_n11_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_5_5_chanX_n3 & track_4_5_chanX_n12 & track_4_6_chanY_n11;
	track_4_5_chanY_n12_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_4_4_chanY_n12 & track_5_4_chanX_n15 & track_4_4_chanX_n4;
	track_4_5_chanY_n13_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_5_5_chanX_n1 & track_4_5_chanX_n14 & track_4_6_chanY_n13;
	track_4_5_chanY_n14_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_4_4_chanY_n14 & track_5_4_chanX_n1 & track_4_4_chanX_n2;
	track_4_5_chanY_n15_driver_mux_fanins <= CLB_5_5_OUT_pin_1 & track_5_5_chanX_n15 & track_4_5_chanX_n0 & track_4_6_chanY_n15;
	track_4_5_chanY_n2_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_4_4_chanY_n2 & track_5_4_chanX_n5 & track_4_4_chanX_n14;
	track_4_5_chanY_n3_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_5_5_chanX_n11 & track_4_5_chanX_n4 & track_4_6_chanY_n3;
	track_4_5_chanY_n4_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_4_4_chanY_n4 & track_5_4_chanX_n7 & track_4_4_chanX_n12;
	track_4_5_chanY_n5_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_5_5_chanX_n9 & track_4_5_chanX_n6 & track_4_6_chanY_n5;
	track_4_5_chanY_n6_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_4_4_chanY_n6 & track_5_4_chanX_n9 & track_4_4_chanX_n10;
	track_4_5_chanY_n7_driver_mux_fanins  <= CLB_4_5_OUT_pin_3 & track_5_5_chanX_n7 & track_4_5_chanX_n8 & track_4_6_chanY_n7;
	track_4_5_chanY_n8_driver_mux_fanins  <= CLB_5_5_OUT_pin_1 & track_4_4_chanY_n8 & track_5_4_chanX_n11 & track_4_4_chanX_n8;
	track_4_5_chanY_n9_driver_mux_fanins  <= CLB_5_5_OUT_pin_1 & track_5_5_chanX_n5 & track_4_5_chanX_n10 & track_4_6_chanY_n9;
	track_4_6_chanX_n0_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_3_6_chanY_n0 & track_3_6_chanX_n0;
	track_4_6_chanX_n1_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_4_6_chanY_n0 & track_5_6_chanX_n1;
	track_4_6_chanX_n10_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_3_6_chanY_n10 & track_3_6_chanX_n10;
	track_4_6_chanX_n11_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_4_6_chanY_n10 & track_5_6_chanX_n11;
	track_4_6_chanX_n12_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_3_6_chanY_n12 & track_3_6_chanX_n12;
	track_4_6_chanX_n13_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_4_6_chanY_n12 & track_5_6_chanX_n13;
	track_4_6_chanX_n14_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_3_6_chanY_n14 & track_3_6_chanX_n14;
	track_4_6_chanX_n15_driver_mux_fanins <= "0" & IO_4_7_OUT_pin_0 & track_4_6_chanY_n14 & track_5_6_chanX_n15;
	track_4_6_chanX_n2_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_3_6_chanY_n2 & track_3_6_chanX_n2;
	track_4_6_chanX_n3_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_4_6_chanY_n2 & track_5_6_chanX_n3;
	track_4_6_chanX_n4_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_3_6_chanY_n4 & track_3_6_chanX_n4;
	track_4_6_chanX_n5_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_4_6_chanY_n4 & track_5_6_chanX_n5;
	track_4_6_chanX_n6_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_3_6_chanY_n6 & track_3_6_chanX_n6;
	track_4_6_chanX_n7_driver_mux_fanins  <= IO_4_7_OUT_pin_1 & CLB_4_6_OUT_pin_2 & track_4_6_chanY_n6 & track_5_6_chanX_n7;
	track_4_6_chanX_n8_driver_mux_fanins  <= "0" & IO_4_7_OUT_pin_0 & track_3_6_chanY_n8 & track_3_6_chanX_n8;
	track_4_6_chanX_n9_driver_mux_fanins  <= "0" & IO_4_7_OUT_pin_0 & track_4_6_chanY_n8 & track_5_6_chanX_n9;
	track_4_6_chanY_n0_driver_mux_fanins  <= CLB_4_6_OUT_pin_3 & track_4_5_chanY_n0 & track_5_5_chanX_n3 & track_4_5_chanX_n0;
	track_4_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_4_6_OUT_pin_3 & track_5_6_chanX_n1 & track_4_6_chanX_n0;
	track_4_6_chanY_n10_driver_mux_fanins <= CLB_5_6_OUT_pin_1 & track_4_5_chanY_n10 & track_5_5_chanX_n13 & track_4_5_chanX_n6;
	track_4_6_chanY_n11_driver_mux_fanins <= "0" & CLB_5_6_OUT_pin_1 & track_5_6_chanX_n5 & track_4_6_chanX_n4;
	track_4_6_chanY_n12_driver_mux_fanins <= CLB_5_6_OUT_pin_1 & track_4_5_chanY_n12 & track_5_5_chanX_n15 & track_4_5_chanX_n4;
	track_4_6_chanY_n13_driver_mux_fanins <= "0" & CLB_5_6_OUT_pin_1 & track_5_6_chanX_n7 & track_4_6_chanX_n6;
	track_4_6_chanY_n14_driver_mux_fanins <= CLB_5_6_OUT_pin_1 & track_4_5_chanY_n14 & track_5_5_chanX_n1 & track_4_5_chanX_n2;
	track_4_6_chanY_n15_driver_mux_fanins <= "0" & CLB_5_6_OUT_pin_1 & track_5_6_chanX_n15 & track_4_6_chanX_n14;
	track_4_6_chanY_n2_driver_mux_fanins  <= CLB_4_6_OUT_pin_3 & track_4_5_chanY_n2 & track_5_5_chanX_n5 & track_4_5_chanX_n14;
	track_4_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_4_6_OUT_pin_3 & track_5_6_chanX_n9 & track_4_6_chanX_n8;
	track_4_6_chanY_n4_driver_mux_fanins  <= CLB_4_6_OUT_pin_3 & track_4_5_chanY_n4 & track_5_5_chanX_n7 & track_4_5_chanX_n12;
	track_4_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_4_6_OUT_pin_3 & track_5_6_chanX_n11 & track_4_6_chanX_n10;
	track_4_6_chanY_n6_driver_mux_fanins  <= CLB_4_6_OUT_pin_3 & track_4_5_chanY_n6 & track_5_5_chanX_n9 & track_4_5_chanX_n10;
	track_4_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_4_6_OUT_pin_3 & track_5_6_chanX_n13 & track_4_6_chanX_n12;
	track_4_6_chanY_n8_driver_mux_fanins  <= CLB_5_6_OUT_pin_1 & track_4_5_chanY_n8 & track_5_5_chanX_n11 & track_4_5_chanX_n8;
	track_4_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_5_6_OUT_pin_1 & track_5_6_chanX_n3 & track_4_6_chanX_n2;
	track_5_0_chanX_n0_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_4_0_chanX_n0 & track_4_1_chanY_n1;
	track_5_0_chanX_n1_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_6_0_chanX_n1 & track_5_1_chanY_n1;
	track_5_0_chanX_n10_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_4_0_chanX_n10 & track_4_1_chanY_n11;
	track_5_0_chanX_n11_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_6_0_chanX_n11 & track_5_1_chanY_n11;
	track_5_0_chanX_n12_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_4_0_chanX_n12 & track_4_1_chanY_n13;
	track_5_0_chanX_n13_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_6_0_chanX_n13 & track_5_1_chanY_n13;
	track_5_0_chanX_n14_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_4_0_chanX_n14 & track_4_1_chanY_n15;
	track_5_0_chanX_n15_driver_mux_fanins <= "0" & IO_5_0_OUT_pin_1 & track_6_0_chanX_n15 & track_5_1_chanY_n15;
	track_5_0_chanX_n2_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_4_0_chanX_n2 & track_4_1_chanY_n3;
	track_5_0_chanX_n3_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_6_0_chanX_n3 & track_5_1_chanY_n3;
	track_5_0_chanX_n4_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_4_0_chanX_n4 & track_4_1_chanY_n5;
	track_5_0_chanX_n5_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_6_0_chanX_n5 & track_5_1_chanY_n5;
	track_5_0_chanX_n6_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_4_0_chanX_n6 & track_4_1_chanY_n7;
	track_5_0_chanX_n7_driver_mux_fanins  <= IO_5_0_OUT_pin_0 & CLB_5_1_OUT_pin_0 & track_6_0_chanX_n7 & track_5_1_chanY_n7;
	track_5_0_chanX_n8_driver_mux_fanins  <= "0" & IO_5_0_OUT_pin_1 & track_4_0_chanX_n8 & track_4_1_chanY_n9;
	track_5_0_chanX_n9_driver_mux_fanins  <= "0" & IO_5_0_OUT_pin_1 & track_6_0_chanX_n9 & track_5_1_chanY_n9;
	track_5_1_chanX_n0_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_4_1_chanY_n12 & track_4_1_chanX_n0 & track_4_2_chanY_n15;
	track_5_1_chanX_n1_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_5_1_chanY_n14 & track_6_1_chanX_n1 & track_5_2_chanY_n1;
	track_5_1_chanX_n10_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_4_1_chanY_n2 & track_4_1_chanX_n10 & track_4_2_chanY_n9;
	track_5_1_chanX_n11_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_5_1_chanY_n8 & track_6_1_chanX_n11 & track_5_2_chanY_n7;
	track_5_1_chanX_n12_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_4_1_chanY_n0 & track_4_1_chanX_n12 & track_4_2_chanY_n11;
	track_5_1_chanX_n13_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_5_1_chanY_n10 & track_6_1_chanX_n13 & track_5_2_chanY_n5;
	track_5_1_chanX_n14_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_4_1_chanY_n14 & track_4_1_chanX_n14 & track_4_2_chanY_n13;
	track_5_1_chanX_n15_driver_mux_fanins <= CLB_5_2_OUT_pin_0 & track_5_1_chanY_n12 & track_6_1_chanX_n15 & track_5_2_chanY_n3;
	track_5_1_chanX_n2_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_4_1_chanY_n10 & track_4_1_chanX_n2 & track_4_2_chanY_n1;
	track_5_1_chanX_n3_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_5_1_chanY_n0 & track_6_1_chanX_n3 & track_5_2_chanY_n15;
	track_5_1_chanX_n4_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_4_1_chanY_n8 & track_4_1_chanX_n4 & track_4_2_chanY_n3;
	track_5_1_chanX_n5_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_5_1_chanY_n2 & track_6_1_chanX_n5 & track_5_2_chanY_n13;
	track_5_1_chanX_n6_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_4_1_chanY_n6 & track_4_1_chanX_n6 & track_4_2_chanY_n5;
	track_5_1_chanX_n7_driver_mux_fanins  <= CLB_5_1_OUT_pin_2 & track_5_1_chanY_n4 & track_6_1_chanX_n7 & track_5_2_chanY_n11;
	track_5_1_chanX_n8_driver_mux_fanins  <= CLB_5_2_OUT_pin_0 & track_4_1_chanY_n4 & track_4_1_chanX_n8 & track_4_2_chanY_n7;
	track_5_1_chanX_n9_driver_mux_fanins  <= CLB_5_2_OUT_pin_0 & track_5_1_chanY_n6 & track_6_1_chanX_n9 & track_5_2_chanY_n9;
	track_5_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_5_1_OUT_pin_3 & track_6_0_chanX_n7 & track_5_0_chanX_n6;
	track_5_1_chanY_n1_driver_mux_fanins  <= CLB_5_1_OUT_pin_3 & track_6_1_chanX_n13 & track_5_1_chanX_n2 & track_5_2_chanY_n1;
	track_5_1_chanY_n10_driver_mux_fanins <= "0" & CLB_6_1_OUT_pin_1 & track_6_0_chanX_n11 & track_5_0_chanX_n10;
	track_5_1_chanY_n11_driver_mux_fanins <= CLB_6_1_OUT_pin_1 & track_6_1_chanX_n3 & track_5_1_chanX_n12 & track_5_2_chanY_n11;
	track_5_1_chanY_n12_driver_mux_fanins <= "0" & CLB_6_1_OUT_pin_1 & track_6_0_chanX_n13 & track_5_0_chanX_n12;
	track_5_1_chanY_n13_driver_mux_fanins <= CLB_6_1_OUT_pin_1 & track_6_1_chanX_n1 & track_5_1_chanX_n14 & track_5_2_chanY_n13;
	track_5_1_chanY_n14_driver_mux_fanins <= "0" & CLB_6_1_OUT_pin_1 & track_6_0_chanX_n15 & track_5_0_chanX_n14;
	track_5_1_chanY_n15_driver_mux_fanins <= CLB_6_1_OUT_pin_1 & track_6_1_chanX_n15 & track_5_1_chanX_n0 & track_5_2_chanY_n15;
	track_5_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_5_1_OUT_pin_3 & track_6_0_chanX_n9 & track_5_0_chanX_n8;
	track_5_1_chanY_n3_driver_mux_fanins  <= CLB_5_1_OUT_pin_3 & track_6_1_chanX_n11 & track_5_1_chanX_n4 & track_5_2_chanY_n3;
	track_5_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_5_1_OUT_pin_3 & track_6_0_chanX_n1 & track_5_0_chanX_n0;
	track_5_1_chanY_n5_driver_mux_fanins  <= CLB_5_1_OUT_pin_3 & track_6_1_chanX_n9 & track_5_1_chanX_n6 & track_5_2_chanY_n5;
	track_5_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_5_1_OUT_pin_3 & track_6_0_chanX_n3 & track_5_0_chanX_n2;
	track_5_1_chanY_n7_driver_mux_fanins  <= CLB_5_1_OUT_pin_3 & track_6_1_chanX_n7 & track_5_1_chanX_n8 & track_5_2_chanY_n7;
	track_5_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_6_1_OUT_pin_1 & track_6_0_chanX_n5 & track_5_0_chanX_n4;
	track_5_1_chanY_n9_driver_mux_fanins  <= CLB_6_1_OUT_pin_1 & track_6_1_chanX_n5 & track_5_1_chanX_n10 & track_5_2_chanY_n9;
	track_5_2_chanX_n0_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_4_2_chanY_n12 & track_4_2_chanX_n0 & track_4_3_chanY_n15;
	track_5_2_chanX_n1_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_5_2_chanY_n14 & track_6_2_chanX_n1 & track_5_3_chanY_n1;
	track_5_2_chanX_n10_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_4_2_chanY_n2 & track_4_2_chanX_n10 & track_4_3_chanY_n9;
	track_5_2_chanX_n11_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_5_2_chanY_n8 & track_6_2_chanX_n11 & track_5_3_chanY_n7;
	track_5_2_chanX_n12_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_4_2_chanY_n0 & track_4_2_chanX_n12 & track_4_3_chanY_n11;
	track_5_2_chanX_n13_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_5_2_chanY_n10 & track_6_2_chanX_n13 & track_5_3_chanY_n5;
	track_5_2_chanX_n14_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_4_2_chanY_n14 & track_4_2_chanX_n14 & track_4_3_chanY_n13;
	track_5_2_chanX_n15_driver_mux_fanins <= CLB_5_3_OUT_pin_0 & track_5_2_chanY_n12 & track_6_2_chanX_n15 & track_5_3_chanY_n3;
	track_5_2_chanX_n2_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_4_2_chanY_n10 & track_4_2_chanX_n2 & track_4_3_chanY_n1;
	track_5_2_chanX_n3_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_5_2_chanY_n0 & track_6_2_chanX_n3 & track_5_3_chanY_n15;
	track_5_2_chanX_n4_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_4_2_chanY_n8 & track_4_2_chanX_n4 & track_4_3_chanY_n3;
	track_5_2_chanX_n5_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_5_2_chanY_n2 & track_6_2_chanX_n5 & track_5_3_chanY_n13;
	track_5_2_chanX_n6_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_4_2_chanY_n6 & track_4_2_chanX_n6 & track_4_3_chanY_n5;
	track_5_2_chanX_n7_driver_mux_fanins  <= CLB_5_2_OUT_pin_2 & track_5_2_chanY_n4 & track_6_2_chanX_n7 & track_5_3_chanY_n11;
	track_5_2_chanX_n8_driver_mux_fanins  <= CLB_5_3_OUT_pin_0 & track_4_2_chanY_n4 & track_4_2_chanX_n8 & track_4_3_chanY_n7;
	track_5_2_chanX_n9_driver_mux_fanins  <= CLB_5_3_OUT_pin_0 & track_5_2_chanY_n6 & track_6_2_chanX_n9 & track_5_3_chanY_n9;
	track_5_2_chanY_n0_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_5_1_chanY_n0 & track_6_1_chanX_n3 & track_5_1_chanX_n0;
	track_5_2_chanY_n1_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_6_2_chanX_n13 & track_5_2_chanX_n2 & track_5_3_chanY_n1;
	track_5_2_chanY_n10_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_5_1_chanY_n10 & track_6_1_chanX_n13 & track_5_1_chanX_n6;
	track_5_2_chanY_n11_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_6_2_chanX_n3 & track_5_2_chanX_n12 & track_5_3_chanY_n11;
	track_5_2_chanY_n12_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_5_1_chanY_n12 & track_6_1_chanX_n15 & track_5_1_chanX_n4;
	track_5_2_chanY_n13_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_6_2_chanX_n1 & track_5_2_chanX_n14 & track_5_3_chanY_n13;
	track_5_2_chanY_n14_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_5_1_chanY_n14 & track_6_1_chanX_n1 & track_5_1_chanX_n2;
	track_5_2_chanY_n15_driver_mux_fanins <= CLB_6_2_OUT_pin_1 & track_6_2_chanX_n15 & track_5_2_chanX_n0 & track_5_3_chanY_n15;
	track_5_2_chanY_n2_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_5_1_chanY_n2 & track_6_1_chanX_n5 & track_5_1_chanX_n14;
	track_5_2_chanY_n3_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_6_2_chanX_n11 & track_5_2_chanX_n4 & track_5_3_chanY_n3;
	track_5_2_chanY_n4_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_5_1_chanY_n4 & track_6_1_chanX_n7 & track_5_1_chanX_n12;
	track_5_2_chanY_n5_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_6_2_chanX_n9 & track_5_2_chanX_n6 & track_5_3_chanY_n5;
	track_5_2_chanY_n6_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_5_1_chanY_n6 & track_6_1_chanX_n9 & track_5_1_chanX_n10;
	track_5_2_chanY_n7_driver_mux_fanins  <= CLB_5_2_OUT_pin_3 & track_6_2_chanX_n7 & track_5_2_chanX_n8 & track_5_3_chanY_n7;
	track_5_2_chanY_n8_driver_mux_fanins  <= CLB_6_2_OUT_pin_1 & track_5_1_chanY_n8 & track_6_1_chanX_n11 & track_5_1_chanX_n8;
	track_5_2_chanY_n9_driver_mux_fanins  <= CLB_6_2_OUT_pin_1 & track_6_2_chanX_n5 & track_5_2_chanX_n10 & track_5_3_chanY_n9;
	track_5_3_chanX_n0_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_4_3_chanY_n12 & track_4_3_chanX_n0 & track_4_4_chanY_n15;
	track_5_3_chanX_n1_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_5_3_chanY_n14 & track_6_3_chanX_n1 & track_5_4_chanY_n1;
	track_5_3_chanX_n10_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_4_3_chanY_n2 & track_4_3_chanX_n10 & track_4_4_chanY_n9;
	track_5_3_chanX_n11_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_5_3_chanY_n8 & track_6_3_chanX_n11 & track_5_4_chanY_n7;
	track_5_3_chanX_n12_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_4_3_chanY_n0 & track_4_3_chanX_n12 & track_4_4_chanY_n11;
	track_5_3_chanX_n13_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_5_3_chanY_n10 & track_6_3_chanX_n13 & track_5_4_chanY_n5;
	track_5_3_chanX_n14_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_4_3_chanY_n14 & track_4_3_chanX_n14 & track_4_4_chanY_n13;
	track_5_3_chanX_n15_driver_mux_fanins <= CLB_5_4_OUT_pin_0 & track_5_3_chanY_n12 & track_6_3_chanX_n15 & track_5_4_chanY_n3;
	track_5_3_chanX_n2_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_4_3_chanY_n10 & track_4_3_chanX_n2 & track_4_4_chanY_n1;
	track_5_3_chanX_n3_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_5_3_chanY_n0 & track_6_3_chanX_n3 & track_5_4_chanY_n15;
	track_5_3_chanX_n4_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_4_3_chanY_n8 & track_4_3_chanX_n4 & track_4_4_chanY_n3;
	track_5_3_chanX_n5_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_5_3_chanY_n2 & track_6_3_chanX_n5 & track_5_4_chanY_n13;
	track_5_3_chanX_n6_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_4_3_chanY_n6 & track_4_3_chanX_n6 & track_4_4_chanY_n5;
	track_5_3_chanX_n7_driver_mux_fanins  <= CLB_5_3_OUT_pin_2 & track_5_3_chanY_n4 & track_6_3_chanX_n7 & track_5_4_chanY_n11;
	track_5_3_chanX_n8_driver_mux_fanins  <= CLB_5_4_OUT_pin_0 & track_4_3_chanY_n4 & track_4_3_chanX_n8 & track_4_4_chanY_n7;
	track_5_3_chanX_n9_driver_mux_fanins  <= CLB_5_4_OUT_pin_0 & track_5_3_chanY_n6 & track_6_3_chanX_n9 & track_5_4_chanY_n9;
	track_5_3_chanY_n0_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_5_2_chanY_n0 & track_6_2_chanX_n3 & track_5_2_chanX_n0;
	track_5_3_chanY_n1_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_6_3_chanX_n13 & track_5_3_chanX_n2 & track_5_4_chanY_n1;
	track_5_3_chanY_n10_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_5_2_chanY_n10 & track_6_2_chanX_n13 & track_5_2_chanX_n6;
	track_5_3_chanY_n11_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_6_3_chanX_n3 & track_5_3_chanX_n12 & track_5_4_chanY_n11;
	track_5_3_chanY_n12_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_5_2_chanY_n12 & track_6_2_chanX_n15 & track_5_2_chanX_n4;
	track_5_3_chanY_n13_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_6_3_chanX_n1 & track_5_3_chanX_n14 & track_5_4_chanY_n13;
	track_5_3_chanY_n14_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_5_2_chanY_n14 & track_6_2_chanX_n1 & track_5_2_chanX_n2;
	track_5_3_chanY_n15_driver_mux_fanins <= CLB_6_3_OUT_pin_1 & track_6_3_chanX_n15 & track_5_3_chanX_n0 & track_5_4_chanY_n15;
	track_5_3_chanY_n2_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_5_2_chanY_n2 & track_6_2_chanX_n5 & track_5_2_chanX_n14;
	track_5_3_chanY_n3_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_6_3_chanX_n11 & track_5_3_chanX_n4 & track_5_4_chanY_n3;
	track_5_3_chanY_n4_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_5_2_chanY_n4 & track_6_2_chanX_n7 & track_5_2_chanX_n12;
	track_5_3_chanY_n5_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_6_3_chanX_n9 & track_5_3_chanX_n6 & track_5_4_chanY_n5;
	track_5_3_chanY_n6_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_5_2_chanY_n6 & track_6_2_chanX_n9 & track_5_2_chanX_n10;
	track_5_3_chanY_n7_driver_mux_fanins  <= CLB_5_3_OUT_pin_3 & track_6_3_chanX_n7 & track_5_3_chanX_n8 & track_5_4_chanY_n7;
	track_5_3_chanY_n8_driver_mux_fanins  <= CLB_6_3_OUT_pin_1 & track_5_2_chanY_n8 & track_6_2_chanX_n11 & track_5_2_chanX_n8;
	track_5_3_chanY_n9_driver_mux_fanins  <= CLB_6_3_OUT_pin_1 & track_6_3_chanX_n5 & track_5_3_chanX_n10 & track_5_4_chanY_n9;
	track_5_4_chanX_n0_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_4_4_chanY_n12 & track_4_4_chanX_n0 & track_4_5_chanY_n15;
	track_5_4_chanX_n1_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_5_4_chanY_n14 & track_6_4_chanX_n1 & track_5_5_chanY_n1;
	track_5_4_chanX_n10_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_4_4_chanY_n2 & track_4_4_chanX_n10 & track_4_5_chanY_n9;
	track_5_4_chanX_n11_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_5_4_chanY_n8 & track_6_4_chanX_n11 & track_5_5_chanY_n7;
	track_5_4_chanX_n12_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_4_4_chanY_n0 & track_4_4_chanX_n12 & track_4_5_chanY_n11;
	track_5_4_chanX_n13_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_5_4_chanY_n10 & track_6_4_chanX_n13 & track_5_5_chanY_n5;
	track_5_4_chanX_n14_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_4_4_chanY_n14 & track_4_4_chanX_n14 & track_4_5_chanY_n13;
	track_5_4_chanX_n15_driver_mux_fanins <= CLB_5_5_OUT_pin_0 & track_5_4_chanY_n12 & track_6_4_chanX_n15 & track_5_5_chanY_n3;
	track_5_4_chanX_n2_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_4_4_chanY_n10 & track_4_4_chanX_n2 & track_4_5_chanY_n1;
	track_5_4_chanX_n3_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_5_4_chanY_n0 & track_6_4_chanX_n3 & track_5_5_chanY_n15;
	track_5_4_chanX_n4_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_4_4_chanY_n8 & track_4_4_chanX_n4 & track_4_5_chanY_n3;
	track_5_4_chanX_n5_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_5_4_chanY_n2 & track_6_4_chanX_n5 & track_5_5_chanY_n13;
	track_5_4_chanX_n6_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_4_4_chanY_n6 & track_4_4_chanX_n6 & track_4_5_chanY_n5;
	track_5_4_chanX_n7_driver_mux_fanins  <= CLB_5_4_OUT_pin_2 & track_5_4_chanY_n4 & track_6_4_chanX_n7 & track_5_5_chanY_n11;
	track_5_4_chanX_n8_driver_mux_fanins  <= CLB_5_5_OUT_pin_0 & track_4_4_chanY_n4 & track_4_4_chanX_n8 & track_4_5_chanY_n7;
	track_5_4_chanX_n9_driver_mux_fanins  <= CLB_5_5_OUT_pin_0 & track_5_4_chanY_n6 & track_6_4_chanX_n9 & track_5_5_chanY_n9;
	track_5_4_chanY_n0_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_5_3_chanY_n0 & track_6_3_chanX_n3 & track_5_3_chanX_n0;
	track_5_4_chanY_n1_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_6_4_chanX_n13 & track_5_4_chanX_n2 & track_5_5_chanY_n1;
	track_5_4_chanY_n10_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_5_3_chanY_n10 & track_6_3_chanX_n13 & track_5_3_chanX_n6;
	track_5_4_chanY_n11_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_6_4_chanX_n3 & track_5_4_chanX_n12 & track_5_5_chanY_n11;
	track_5_4_chanY_n12_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_5_3_chanY_n12 & track_6_3_chanX_n15 & track_5_3_chanX_n4;
	track_5_4_chanY_n13_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_6_4_chanX_n1 & track_5_4_chanX_n14 & track_5_5_chanY_n13;
	track_5_4_chanY_n14_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_5_3_chanY_n14 & track_6_3_chanX_n1 & track_5_3_chanX_n2;
	track_5_4_chanY_n15_driver_mux_fanins <= CLB_6_4_OUT_pin_1 & track_6_4_chanX_n15 & track_5_4_chanX_n0 & track_5_5_chanY_n15;
	track_5_4_chanY_n2_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_5_3_chanY_n2 & track_6_3_chanX_n5 & track_5_3_chanX_n14;
	track_5_4_chanY_n3_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_6_4_chanX_n11 & track_5_4_chanX_n4 & track_5_5_chanY_n3;
	track_5_4_chanY_n4_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_5_3_chanY_n4 & track_6_3_chanX_n7 & track_5_3_chanX_n12;
	track_5_4_chanY_n5_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_6_4_chanX_n9 & track_5_4_chanX_n6 & track_5_5_chanY_n5;
	track_5_4_chanY_n6_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_5_3_chanY_n6 & track_6_3_chanX_n9 & track_5_3_chanX_n10;
	track_5_4_chanY_n7_driver_mux_fanins  <= CLB_5_4_OUT_pin_3 & track_6_4_chanX_n7 & track_5_4_chanX_n8 & track_5_5_chanY_n7;
	track_5_4_chanY_n8_driver_mux_fanins  <= CLB_6_4_OUT_pin_1 & track_5_3_chanY_n8 & track_6_3_chanX_n11 & track_5_3_chanX_n8;
	track_5_4_chanY_n9_driver_mux_fanins  <= CLB_6_4_OUT_pin_1 & track_6_4_chanX_n5 & track_5_4_chanX_n10 & track_5_5_chanY_n9;
	track_5_5_chanX_n0_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_4_5_chanY_n12 & track_4_5_chanX_n0 & track_4_6_chanY_n15;
	track_5_5_chanX_n1_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_5_5_chanY_n14 & track_6_5_chanX_n1 & track_5_6_chanY_n1;
	track_5_5_chanX_n10_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_4_5_chanY_n2 & track_4_5_chanX_n10 & track_4_6_chanY_n9;
	track_5_5_chanX_n11_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_5_5_chanY_n8 & track_6_5_chanX_n11 & track_5_6_chanY_n7;
	track_5_5_chanX_n12_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_4_5_chanY_n0 & track_4_5_chanX_n12 & track_4_6_chanY_n11;
	track_5_5_chanX_n13_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_5_5_chanY_n10 & track_6_5_chanX_n13 & track_5_6_chanY_n5;
	track_5_5_chanX_n14_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_4_5_chanY_n14 & track_4_5_chanX_n14 & track_4_6_chanY_n13;
	track_5_5_chanX_n15_driver_mux_fanins <= CLB_5_6_OUT_pin_0 & track_5_5_chanY_n12 & track_6_5_chanX_n15 & track_5_6_chanY_n3;
	track_5_5_chanX_n2_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_4_5_chanY_n10 & track_4_5_chanX_n2 & track_4_6_chanY_n1;
	track_5_5_chanX_n3_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_5_5_chanY_n0 & track_6_5_chanX_n3 & track_5_6_chanY_n15;
	track_5_5_chanX_n4_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_4_5_chanY_n8 & track_4_5_chanX_n4 & track_4_6_chanY_n3;
	track_5_5_chanX_n5_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_5_5_chanY_n2 & track_6_5_chanX_n5 & track_5_6_chanY_n13;
	track_5_5_chanX_n6_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_4_5_chanY_n6 & track_4_5_chanX_n6 & track_4_6_chanY_n5;
	track_5_5_chanX_n7_driver_mux_fanins  <= CLB_5_5_OUT_pin_2 & track_5_5_chanY_n4 & track_6_5_chanX_n7 & track_5_6_chanY_n11;
	track_5_5_chanX_n8_driver_mux_fanins  <= CLB_5_6_OUT_pin_0 & track_4_5_chanY_n4 & track_4_5_chanX_n8 & track_4_6_chanY_n7;
	track_5_5_chanX_n9_driver_mux_fanins  <= CLB_5_6_OUT_pin_0 & track_5_5_chanY_n6 & track_6_5_chanX_n9 & track_5_6_chanY_n9;
	track_5_5_chanY_n0_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_5_4_chanY_n0 & track_6_4_chanX_n3 & track_5_4_chanX_n0;
	track_5_5_chanY_n1_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_6_5_chanX_n13 & track_5_5_chanX_n2 & track_5_6_chanY_n1;
	track_5_5_chanY_n10_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_5_4_chanY_n10 & track_6_4_chanX_n13 & track_5_4_chanX_n6;
	track_5_5_chanY_n11_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_6_5_chanX_n3 & track_5_5_chanX_n12 & track_5_6_chanY_n11;
	track_5_5_chanY_n12_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_5_4_chanY_n12 & track_6_4_chanX_n15 & track_5_4_chanX_n4;
	track_5_5_chanY_n13_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_6_5_chanX_n1 & track_5_5_chanX_n14 & track_5_6_chanY_n13;
	track_5_5_chanY_n14_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_5_4_chanY_n14 & track_6_4_chanX_n1 & track_5_4_chanX_n2;
	track_5_5_chanY_n15_driver_mux_fanins <= CLB_6_5_OUT_pin_1 & track_6_5_chanX_n15 & track_5_5_chanX_n0 & track_5_6_chanY_n15;
	track_5_5_chanY_n2_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_5_4_chanY_n2 & track_6_4_chanX_n5 & track_5_4_chanX_n14;
	track_5_5_chanY_n3_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_6_5_chanX_n11 & track_5_5_chanX_n4 & track_5_6_chanY_n3;
	track_5_5_chanY_n4_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_5_4_chanY_n4 & track_6_4_chanX_n7 & track_5_4_chanX_n12;
	track_5_5_chanY_n5_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_6_5_chanX_n9 & track_5_5_chanX_n6 & track_5_6_chanY_n5;
	track_5_5_chanY_n6_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_5_4_chanY_n6 & track_6_4_chanX_n9 & track_5_4_chanX_n10;
	track_5_5_chanY_n7_driver_mux_fanins  <= CLB_5_5_OUT_pin_3 & track_6_5_chanX_n7 & track_5_5_chanX_n8 & track_5_6_chanY_n7;
	track_5_5_chanY_n8_driver_mux_fanins  <= CLB_6_5_OUT_pin_1 & track_5_4_chanY_n8 & track_6_4_chanX_n11 & track_5_4_chanX_n8;
	track_5_5_chanY_n9_driver_mux_fanins  <= CLB_6_5_OUT_pin_1 & track_6_5_chanX_n5 & track_5_5_chanX_n10 & track_5_6_chanY_n9;
	track_5_6_chanX_n0_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_4_6_chanY_n0 & track_4_6_chanX_n0;
	track_5_6_chanX_n1_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_5_6_chanY_n0 & track_6_6_chanX_n1;
	track_5_6_chanX_n10_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_4_6_chanY_n10 & track_4_6_chanX_n10;
	track_5_6_chanX_n11_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_5_6_chanY_n10 & track_6_6_chanX_n11;
	track_5_6_chanX_n12_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_4_6_chanY_n12 & track_4_6_chanX_n12;
	track_5_6_chanX_n13_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_5_6_chanY_n12 & track_6_6_chanX_n13;
	track_5_6_chanX_n14_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_4_6_chanY_n14 & track_4_6_chanX_n14;
	track_5_6_chanX_n15_driver_mux_fanins <= "0" & IO_5_7_OUT_pin_0 & track_5_6_chanY_n14 & track_6_6_chanX_n15;
	track_5_6_chanX_n2_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_4_6_chanY_n2 & track_4_6_chanX_n2;
	track_5_6_chanX_n3_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_5_6_chanY_n2 & track_6_6_chanX_n3;
	track_5_6_chanX_n4_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_4_6_chanY_n4 & track_4_6_chanX_n4;
	track_5_6_chanX_n5_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_5_6_chanY_n4 & track_6_6_chanX_n5;
	track_5_6_chanX_n6_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_4_6_chanY_n6 & track_4_6_chanX_n6;
	track_5_6_chanX_n7_driver_mux_fanins  <= IO_5_7_OUT_pin_1 & CLB_5_6_OUT_pin_2 & track_5_6_chanY_n6 & track_6_6_chanX_n7;
	track_5_6_chanX_n8_driver_mux_fanins  <= "0" & IO_5_7_OUT_pin_0 & track_4_6_chanY_n8 & track_4_6_chanX_n8;
	track_5_6_chanX_n9_driver_mux_fanins  <= "0" & IO_5_7_OUT_pin_0 & track_5_6_chanY_n8 & track_6_6_chanX_n9;
	track_5_6_chanY_n0_driver_mux_fanins  <= CLB_5_6_OUT_pin_3 & track_5_5_chanY_n0 & track_6_5_chanX_n3 & track_5_5_chanX_n0;
	track_5_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_5_6_OUT_pin_3 & track_6_6_chanX_n1 & track_5_6_chanX_n0;
	track_5_6_chanY_n10_driver_mux_fanins <= CLB_6_6_OUT_pin_1 & track_5_5_chanY_n10 & track_6_5_chanX_n13 & track_5_5_chanX_n6;
	track_5_6_chanY_n11_driver_mux_fanins <= "0" & CLB_6_6_OUT_pin_1 & track_6_6_chanX_n5 & track_5_6_chanX_n4;
	track_5_6_chanY_n12_driver_mux_fanins <= CLB_6_6_OUT_pin_1 & track_5_5_chanY_n12 & track_6_5_chanX_n15 & track_5_5_chanX_n4;
	track_5_6_chanY_n13_driver_mux_fanins <= "0" & CLB_6_6_OUT_pin_1 & track_6_6_chanX_n7 & track_5_6_chanX_n6;
	track_5_6_chanY_n14_driver_mux_fanins <= CLB_6_6_OUT_pin_1 & track_5_5_chanY_n14 & track_6_5_chanX_n1 & track_5_5_chanX_n2;
	track_5_6_chanY_n15_driver_mux_fanins <= "0" & CLB_6_6_OUT_pin_1 & track_6_6_chanX_n15 & track_5_6_chanX_n14;
	track_5_6_chanY_n2_driver_mux_fanins  <= CLB_5_6_OUT_pin_3 & track_5_5_chanY_n2 & track_6_5_chanX_n5 & track_5_5_chanX_n14;
	track_5_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_5_6_OUT_pin_3 & track_6_6_chanX_n9 & track_5_6_chanX_n8;
	track_5_6_chanY_n4_driver_mux_fanins  <= CLB_5_6_OUT_pin_3 & track_5_5_chanY_n4 & track_6_5_chanX_n7 & track_5_5_chanX_n12;
	track_5_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_5_6_OUT_pin_3 & track_6_6_chanX_n11 & track_5_6_chanX_n10;
	track_5_6_chanY_n6_driver_mux_fanins  <= CLB_5_6_OUT_pin_3 & track_5_5_chanY_n6 & track_6_5_chanX_n9 & track_5_5_chanX_n10;
	track_5_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_5_6_OUT_pin_3 & track_6_6_chanX_n13 & track_5_6_chanX_n12;
	track_5_6_chanY_n8_driver_mux_fanins  <= CLB_6_6_OUT_pin_1 & track_5_5_chanY_n8 & track_6_5_chanX_n11 & track_5_5_chanX_n8;
	track_5_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_6_6_OUT_pin_1 & track_6_6_chanX_n3 & track_5_6_chanX_n2;
	track_6_0_chanX_n0_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_5_0_chanX_n0 & track_5_1_chanY_n1;
	track_6_0_chanX_n1_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_7_0_chanX_n1 & track_6_1_chanY_n1;
	track_6_0_chanX_n10_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_5_0_chanX_n10 & track_5_1_chanY_n11;
	track_6_0_chanX_n11_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_7_0_chanX_n11 & track_6_1_chanY_n11;
	track_6_0_chanX_n12_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_5_0_chanX_n12 & track_5_1_chanY_n13;
	track_6_0_chanX_n13_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_7_0_chanX_n13 & track_6_1_chanY_n13;
	track_6_0_chanX_n14_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_5_0_chanX_n14 & track_5_1_chanY_n15;
	track_6_0_chanX_n15_driver_mux_fanins <= "0" & IO_6_0_OUT_pin_1 & track_7_0_chanX_n15 & track_6_1_chanY_n15;
	track_6_0_chanX_n2_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_5_0_chanX_n2 & track_5_1_chanY_n3;
	track_6_0_chanX_n3_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_7_0_chanX_n3 & track_6_1_chanY_n3;
	track_6_0_chanX_n4_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_5_0_chanX_n4 & track_5_1_chanY_n5;
	track_6_0_chanX_n5_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_7_0_chanX_n5 & track_6_1_chanY_n5;
	track_6_0_chanX_n6_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_5_0_chanX_n6 & track_5_1_chanY_n7;
	track_6_0_chanX_n7_driver_mux_fanins  <= IO_6_0_OUT_pin_0 & CLB_6_1_OUT_pin_0 & track_7_0_chanX_n7 & track_6_1_chanY_n7;
	track_6_0_chanX_n8_driver_mux_fanins  <= "0" & IO_6_0_OUT_pin_1 & track_5_0_chanX_n8 & track_5_1_chanY_n9;
	track_6_0_chanX_n9_driver_mux_fanins  <= "0" & IO_6_0_OUT_pin_1 & track_7_0_chanX_n9 & track_6_1_chanY_n9;
	track_6_1_chanX_n0_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_5_1_chanY_n12 & track_5_1_chanX_n0 & track_5_2_chanY_n15;
	track_6_1_chanX_n1_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_6_1_chanY_n14 & track_7_1_chanX_n1 & track_6_2_chanY_n1;
	track_6_1_chanX_n10_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_5_1_chanY_n2 & track_5_1_chanX_n10 & track_5_2_chanY_n9;
	track_6_1_chanX_n11_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_6_1_chanY_n8 & track_7_1_chanX_n11 & track_6_2_chanY_n7;
	track_6_1_chanX_n12_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_5_1_chanY_n0 & track_5_1_chanX_n12 & track_5_2_chanY_n11;
	track_6_1_chanX_n13_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_6_1_chanY_n10 & track_7_1_chanX_n13 & track_6_2_chanY_n5;
	track_6_1_chanX_n14_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_5_1_chanY_n14 & track_5_1_chanX_n14 & track_5_2_chanY_n13;
	track_6_1_chanX_n15_driver_mux_fanins <= CLB_6_2_OUT_pin_0 & track_6_1_chanY_n12 & track_7_1_chanX_n15 & track_6_2_chanY_n3;
	track_6_1_chanX_n2_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_5_1_chanY_n10 & track_5_1_chanX_n2 & track_5_2_chanY_n1;
	track_6_1_chanX_n3_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_6_1_chanY_n0 & track_7_1_chanX_n3 & track_6_2_chanY_n15;
	track_6_1_chanX_n4_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_5_1_chanY_n8 & track_5_1_chanX_n4 & track_5_2_chanY_n3;
	track_6_1_chanX_n5_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_6_1_chanY_n2 & track_7_1_chanX_n5 & track_6_2_chanY_n13;
	track_6_1_chanX_n6_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_5_1_chanY_n6 & track_5_1_chanX_n6 & track_5_2_chanY_n5;
	track_6_1_chanX_n7_driver_mux_fanins  <= CLB_6_1_OUT_pin_2 & track_6_1_chanY_n4 & track_7_1_chanX_n7 & track_6_2_chanY_n11;
	track_6_1_chanX_n8_driver_mux_fanins  <= CLB_6_2_OUT_pin_0 & track_5_1_chanY_n4 & track_5_1_chanX_n8 & track_5_2_chanY_n7;
	track_6_1_chanX_n9_driver_mux_fanins  <= CLB_6_2_OUT_pin_0 & track_6_1_chanY_n6 & track_7_1_chanX_n9 & track_6_2_chanY_n9;
	track_6_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_6_1_OUT_pin_3 & track_7_0_chanX_n7 & track_6_0_chanX_n6;
	track_6_1_chanY_n1_driver_mux_fanins  <= CLB_6_1_OUT_pin_3 & track_7_1_chanX_n13 & track_6_1_chanX_n2 & track_6_2_chanY_n1;
	track_6_1_chanY_n10_driver_mux_fanins <= "0" & CLB_7_1_OUT_pin_1 & track_7_0_chanX_n11 & track_6_0_chanX_n10;
	track_6_1_chanY_n11_driver_mux_fanins <= CLB_7_1_OUT_pin_1 & track_7_1_chanX_n3 & track_6_1_chanX_n12 & track_6_2_chanY_n11;
	track_6_1_chanY_n12_driver_mux_fanins <= "0" & CLB_7_1_OUT_pin_1 & track_7_0_chanX_n13 & track_6_0_chanX_n12;
	track_6_1_chanY_n13_driver_mux_fanins <= CLB_7_1_OUT_pin_1 & track_7_1_chanX_n1 & track_6_1_chanX_n14 & track_6_2_chanY_n13;
	track_6_1_chanY_n14_driver_mux_fanins <= "0" & CLB_7_1_OUT_pin_1 & track_7_0_chanX_n15 & track_6_0_chanX_n14;
	track_6_1_chanY_n15_driver_mux_fanins <= CLB_7_1_OUT_pin_1 & track_7_1_chanX_n15 & track_6_1_chanX_n0 & track_6_2_chanY_n15;
	track_6_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_6_1_OUT_pin_3 & track_7_0_chanX_n9 & track_6_0_chanX_n8;
	track_6_1_chanY_n3_driver_mux_fanins  <= CLB_6_1_OUT_pin_3 & track_7_1_chanX_n11 & track_6_1_chanX_n4 & track_6_2_chanY_n3;
	track_6_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_6_1_OUT_pin_3 & track_7_0_chanX_n1 & track_6_0_chanX_n0;
	track_6_1_chanY_n5_driver_mux_fanins  <= CLB_6_1_OUT_pin_3 & track_7_1_chanX_n9 & track_6_1_chanX_n6 & track_6_2_chanY_n5;
	track_6_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_6_1_OUT_pin_3 & track_7_0_chanX_n3 & track_6_0_chanX_n2;
	track_6_1_chanY_n7_driver_mux_fanins  <= CLB_6_1_OUT_pin_3 & track_7_1_chanX_n7 & track_6_1_chanX_n8 & track_6_2_chanY_n7;
	track_6_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_7_1_OUT_pin_1 & track_7_0_chanX_n5 & track_6_0_chanX_n4;
	track_6_1_chanY_n9_driver_mux_fanins  <= CLB_7_1_OUT_pin_1 & track_7_1_chanX_n5 & track_6_1_chanX_n10 & track_6_2_chanY_n9;
	track_6_2_chanX_n0_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_5_2_chanY_n12 & track_5_2_chanX_n0 & track_5_3_chanY_n15;
	track_6_2_chanX_n1_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_6_2_chanY_n14 & track_7_2_chanX_n1 & track_6_3_chanY_n1;
	track_6_2_chanX_n10_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_5_2_chanY_n2 & track_5_2_chanX_n10 & track_5_3_chanY_n9;
	track_6_2_chanX_n11_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_6_2_chanY_n8 & track_7_2_chanX_n11 & track_6_3_chanY_n7;
	track_6_2_chanX_n12_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_5_2_chanY_n0 & track_5_2_chanX_n12 & track_5_3_chanY_n11;
	track_6_2_chanX_n13_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_6_2_chanY_n10 & track_7_2_chanX_n13 & track_6_3_chanY_n5;
	track_6_2_chanX_n14_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_5_2_chanY_n14 & track_5_2_chanX_n14 & track_5_3_chanY_n13;
	track_6_2_chanX_n15_driver_mux_fanins <= CLB_6_3_OUT_pin_0 & track_6_2_chanY_n12 & track_7_2_chanX_n15 & track_6_3_chanY_n3;
	track_6_2_chanX_n2_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_5_2_chanY_n10 & track_5_2_chanX_n2 & track_5_3_chanY_n1;
	track_6_2_chanX_n3_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_6_2_chanY_n0 & track_7_2_chanX_n3 & track_6_3_chanY_n15;
	track_6_2_chanX_n4_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_5_2_chanY_n8 & track_5_2_chanX_n4 & track_5_3_chanY_n3;
	track_6_2_chanX_n5_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_6_2_chanY_n2 & track_7_2_chanX_n5 & track_6_3_chanY_n13;
	track_6_2_chanX_n6_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_5_2_chanY_n6 & track_5_2_chanX_n6 & track_5_3_chanY_n5;
	track_6_2_chanX_n7_driver_mux_fanins  <= CLB_6_2_OUT_pin_2 & track_6_2_chanY_n4 & track_7_2_chanX_n7 & track_6_3_chanY_n11;
	track_6_2_chanX_n8_driver_mux_fanins  <= CLB_6_3_OUT_pin_0 & track_5_2_chanY_n4 & track_5_2_chanX_n8 & track_5_3_chanY_n7;
	track_6_2_chanX_n9_driver_mux_fanins  <= CLB_6_3_OUT_pin_0 & track_6_2_chanY_n6 & track_7_2_chanX_n9 & track_6_3_chanY_n9;
	track_6_2_chanY_n0_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_6_1_chanY_n0 & track_7_1_chanX_n3 & track_6_1_chanX_n0;
	track_6_2_chanY_n1_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_7_2_chanX_n13 & track_6_2_chanX_n2 & track_6_3_chanY_n1;
	track_6_2_chanY_n10_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_6_1_chanY_n10 & track_7_1_chanX_n13 & track_6_1_chanX_n6;
	track_6_2_chanY_n11_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_7_2_chanX_n3 & track_6_2_chanX_n12 & track_6_3_chanY_n11;
	track_6_2_chanY_n12_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_6_1_chanY_n12 & track_7_1_chanX_n15 & track_6_1_chanX_n4;
	track_6_2_chanY_n13_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_7_2_chanX_n1 & track_6_2_chanX_n14 & track_6_3_chanY_n13;
	track_6_2_chanY_n14_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_6_1_chanY_n14 & track_7_1_chanX_n1 & track_6_1_chanX_n2;
	track_6_2_chanY_n15_driver_mux_fanins <= CLB_7_2_OUT_pin_1 & track_7_2_chanX_n15 & track_6_2_chanX_n0 & track_6_3_chanY_n15;
	track_6_2_chanY_n2_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_6_1_chanY_n2 & track_7_1_chanX_n5 & track_6_1_chanX_n14;
	track_6_2_chanY_n3_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_7_2_chanX_n11 & track_6_2_chanX_n4 & track_6_3_chanY_n3;
	track_6_2_chanY_n4_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_6_1_chanY_n4 & track_7_1_chanX_n7 & track_6_1_chanX_n12;
	track_6_2_chanY_n5_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_7_2_chanX_n9 & track_6_2_chanX_n6 & track_6_3_chanY_n5;
	track_6_2_chanY_n6_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_6_1_chanY_n6 & track_7_1_chanX_n9 & track_6_1_chanX_n10;
	track_6_2_chanY_n7_driver_mux_fanins  <= CLB_6_2_OUT_pin_3 & track_7_2_chanX_n7 & track_6_2_chanX_n8 & track_6_3_chanY_n7;
	track_6_2_chanY_n8_driver_mux_fanins  <= CLB_7_2_OUT_pin_1 & track_6_1_chanY_n8 & track_7_1_chanX_n11 & track_6_1_chanX_n8;
	track_6_2_chanY_n9_driver_mux_fanins  <= CLB_7_2_OUT_pin_1 & track_7_2_chanX_n5 & track_6_2_chanX_n10 & track_6_3_chanY_n9;
	track_6_3_chanX_n0_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_5_3_chanY_n12 & track_5_3_chanX_n0 & track_5_4_chanY_n15;
	track_6_3_chanX_n1_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_6_3_chanY_n14 & track_7_3_chanX_n1 & track_6_4_chanY_n1;
	track_6_3_chanX_n10_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_5_3_chanY_n2 & track_5_3_chanX_n10 & track_5_4_chanY_n9;
	track_6_3_chanX_n11_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_6_3_chanY_n8 & track_7_3_chanX_n11 & track_6_4_chanY_n7;
	track_6_3_chanX_n12_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_5_3_chanY_n0 & track_5_3_chanX_n12 & track_5_4_chanY_n11;
	track_6_3_chanX_n13_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_6_3_chanY_n10 & track_7_3_chanX_n13 & track_6_4_chanY_n5;
	track_6_3_chanX_n14_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_5_3_chanY_n14 & track_5_3_chanX_n14 & track_5_4_chanY_n13;
	track_6_3_chanX_n15_driver_mux_fanins <= CLB_6_4_OUT_pin_0 & track_6_3_chanY_n12 & track_7_3_chanX_n15 & track_6_4_chanY_n3;
	track_6_3_chanX_n2_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_5_3_chanY_n10 & track_5_3_chanX_n2 & track_5_4_chanY_n1;
	track_6_3_chanX_n3_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_6_3_chanY_n0 & track_7_3_chanX_n3 & track_6_4_chanY_n15;
	track_6_3_chanX_n4_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_5_3_chanY_n8 & track_5_3_chanX_n4 & track_5_4_chanY_n3;
	track_6_3_chanX_n5_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_6_3_chanY_n2 & track_7_3_chanX_n5 & track_6_4_chanY_n13;
	track_6_3_chanX_n6_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_5_3_chanY_n6 & track_5_3_chanX_n6 & track_5_4_chanY_n5;
	track_6_3_chanX_n7_driver_mux_fanins  <= CLB_6_3_OUT_pin_2 & track_6_3_chanY_n4 & track_7_3_chanX_n7 & track_6_4_chanY_n11;
	track_6_3_chanX_n8_driver_mux_fanins  <= CLB_6_4_OUT_pin_0 & track_5_3_chanY_n4 & track_5_3_chanX_n8 & track_5_4_chanY_n7;
	track_6_3_chanX_n9_driver_mux_fanins  <= CLB_6_4_OUT_pin_0 & track_6_3_chanY_n6 & track_7_3_chanX_n9 & track_6_4_chanY_n9;
	track_6_3_chanY_n0_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_6_2_chanY_n0 & track_7_2_chanX_n3 & track_6_2_chanX_n0;
	track_6_3_chanY_n1_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_7_3_chanX_n13 & track_6_3_chanX_n2 & track_6_4_chanY_n1;
	track_6_3_chanY_n10_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_6_2_chanY_n10 & track_7_2_chanX_n13 & track_6_2_chanX_n6;
	track_6_3_chanY_n11_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_7_3_chanX_n3 & track_6_3_chanX_n12 & track_6_4_chanY_n11;
	track_6_3_chanY_n12_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_6_2_chanY_n12 & track_7_2_chanX_n15 & track_6_2_chanX_n4;
	track_6_3_chanY_n13_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_7_3_chanX_n1 & track_6_3_chanX_n14 & track_6_4_chanY_n13;
	track_6_3_chanY_n14_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_6_2_chanY_n14 & track_7_2_chanX_n1 & track_6_2_chanX_n2;
	track_6_3_chanY_n15_driver_mux_fanins <= CLB_7_3_OUT_pin_1 & track_7_3_chanX_n15 & track_6_3_chanX_n0 & track_6_4_chanY_n15;
	track_6_3_chanY_n2_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_6_2_chanY_n2 & track_7_2_chanX_n5 & track_6_2_chanX_n14;
	track_6_3_chanY_n3_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_7_3_chanX_n11 & track_6_3_chanX_n4 & track_6_4_chanY_n3;
	track_6_3_chanY_n4_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_6_2_chanY_n4 & track_7_2_chanX_n7 & track_6_2_chanX_n12;
	track_6_3_chanY_n5_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_7_3_chanX_n9 & track_6_3_chanX_n6 & track_6_4_chanY_n5;
	track_6_3_chanY_n6_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_6_2_chanY_n6 & track_7_2_chanX_n9 & track_6_2_chanX_n10;
	track_6_3_chanY_n7_driver_mux_fanins  <= CLB_6_3_OUT_pin_3 & track_7_3_chanX_n7 & track_6_3_chanX_n8 & track_6_4_chanY_n7;
	track_6_3_chanY_n8_driver_mux_fanins  <= CLB_7_3_OUT_pin_1 & track_6_2_chanY_n8 & track_7_2_chanX_n11 & track_6_2_chanX_n8;
	track_6_3_chanY_n9_driver_mux_fanins  <= CLB_7_3_OUT_pin_1 & track_7_3_chanX_n5 & track_6_3_chanX_n10 & track_6_4_chanY_n9;
	track_6_4_chanX_n0_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_5_4_chanY_n12 & track_5_4_chanX_n0 & track_5_5_chanY_n15;
	track_6_4_chanX_n1_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_6_4_chanY_n14 & track_7_4_chanX_n1 & track_6_5_chanY_n1;
	track_6_4_chanX_n10_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_5_4_chanY_n2 & track_5_4_chanX_n10 & track_5_5_chanY_n9;
	track_6_4_chanX_n11_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_6_4_chanY_n8 & track_7_4_chanX_n11 & track_6_5_chanY_n7;
	track_6_4_chanX_n12_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_5_4_chanY_n0 & track_5_4_chanX_n12 & track_5_5_chanY_n11;
	track_6_4_chanX_n13_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_6_4_chanY_n10 & track_7_4_chanX_n13 & track_6_5_chanY_n5;
	track_6_4_chanX_n14_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_5_4_chanY_n14 & track_5_4_chanX_n14 & track_5_5_chanY_n13;
	track_6_4_chanX_n15_driver_mux_fanins <= CLB_6_5_OUT_pin_0 & track_6_4_chanY_n12 & track_7_4_chanX_n15 & track_6_5_chanY_n3;
	track_6_4_chanX_n2_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_5_4_chanY_n10 & track_5_4_chanX_n2 & track_5_5_chanY_n1;
	track_6_4_chanX_n3_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_6_4_chanY_n0 & track_7_4_chanX_n3 & track_6_5_chanY_n15;
	track_6_4_chanX_n4_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_5_4_chanY_n8 & track_5_4_chanX_n4 & track_5_5_chanY_n3;
	track_6_4_chanX_n5_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_6_4_chanY_n2 & track_7_4_chanX_n5 & track_6_5_chanY_n13;
	track_6_4_chanX_n6_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_5_4_chanY_n6 & track_5_4_chanX_n6 & track_5_5_chanY_n5;
	track_6_4_chanX_n7_driver_mux_fanins  <= CLB_6_4_OUT_pin_2 & track_6_4_chanY_n4 & track_7_4_chanX_n7 & track_6_5_chanY_n11;
	track_6_4_chanX_n8_driver_mux_fanins  <= CLB_6_5_OUT_pin_0 & track_5_4_chanY_n4 & track_5_4_chanX_n8 & track_5_5_chanY_n7;
	track_6_4_chanX_n9_driver_mux_fanins  <= CLB_6_5_OUT_pin_0 & track_6_4_chanY_n6 & track_7_4_chanX_n9 & track_6_5_chanY_n9;
	track_6_4_chanY_n0_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_6_3_chanY_n0 & track_7_3_chanX_n3 & track_6_3_chanX_n0;
	track_6_4_chanY_n1_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_7_4_chanX_n13 & track_6_4_chanX_n2 & track_6_5_chanY_n1;
	track_6_4_chanY_n10_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_6_3_chanY_n10 & track_7_3_chanX_n13 & track_6_3_chanX_n6;
	track_6_4_chanY_n11_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_7_4_chanX_n3 & track_6_4_chanX_n12 & track_6_5_chanY_n11;
	track_6_4_chanY_n12_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_6_3_chanY_n12 & track_7_3_chanX_n15 & track_6_3_chanX_n4;
	track_6_4_chanY_n13_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_7_4_chanX_n1 & track_6_4_chanX_n14 & track_6_5_chanY_n13;
	track_6_4_chanY_n14_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_6_3_chanY_n14 & track_7_3_chanX_n1 & track_6_3_chanX_n2;
	track_6_4_chanY_n15_driver_mux_fanins <= CLB_7_4_OUT_pin_1 & track_7_4_chanX_n15 & track_6_4_chanX_n0 & track_6_5_chanY_n15;
	track_6_4_chanY_n2_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_6_3_chanY_n2 & track_7_3_chanX_n5 & track_6_3_chanX_n14;
	track_6_4_chanY_n3_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_7_4_chanX_n11 & track_6_4_chanX_n4 & track_6_5_chanY_n3;
	track_6_4_chanY_n4_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_6_3_chanY_n4 & track_7_3_chanX_n7 & track_6_3_chanX_n12;
	track_6_4_chanY_n5_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_7_4_chanX_n9 & track_6_4_chanX_n6 & track_6_5_chanY_n5;
	track_6_4_chanY_n6_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_6_3_chanY_n6 & track_7_3_chanX_n9 & track_6_3_chanX_n10;
	track_6_4_chanY_n7_driver_mux_fanins  <= CLB_6_4_OUT_pin_3 & track_7_4_chanX_n7 & track_6_4_chanX_n8 & track_6_5_chanY_n7;
	track_6_4_chanY_n8_driver_mux_fanins  <= CLB_7_4_OUT_pin_1 & track_6_3_chanY_n8 & track_7_3_chanX_n11 & track_6_3_chanX_n8;
	track_6_4_chanY_n9_driver_mux_fanins  <= CLB_7_4_OUT_pin_1 & track_7_4_chanX_n5 & track_6_4_chanX_n10 & track_6_5_chanY_n9;
	track_6_5_chanX_n0_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_5_5_chanY_n12 & track_5_5_chanX_n0 & track_5_6_chanY_n15;
	track_6_5_chanX_n1_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_6_5_chanY_n14 & track_7_5_chanX_n1 & track_6_6_chanY_n1;
	track_6_5_chanX_n10_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_5_5_chanY_n2 & track_5_5_chanX_n10 & track_5_6_chanY_n9;
	track_6_5_chanX_n11_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_6_5_chanY_n8 & track_7_5_chanX_n11 & track_6_6_chanY_n7;
	track_6_5_chanX_n12_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_5_5_chanY_n0 & track_5_5_chanX_n12 & track_5_6_chanY_n11;
	track_6_5_chanX_n13_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_6_5_chanY_n10 & track_7_5_chanX_n13 & track_6_6_chanY_n5;
	track_6_5_chanX_n14_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_5_5_chanY_n14 & track_5_5_chanX_n14 & track_5_6_chanY_n13;
	track_6_5_chanX_n15_driver_mux_fanins <= CLB_6_6_OUT_pin_0 & track_6_5_chanY_n12 & track_7_5_chanX_n15 & track_6_6_chanY_n3;
	track_6_5_chanX_n2_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_5_5_chanY_n10 & track_5_5_chanX_n2 & track_5_6_chanY_n1;
	track_6_5_chanX_n3_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_6_5_chanY_n0 & track_7_5_chanX_n3 & track_6_6_chanY_n15;
	track_6_5_chanX_n4_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_5_5_chanY_n8 & track_5_5_chanX_n4 & track_5_6_chanY_n3;
	track_6_5_chanX_n5_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_6_5_chanY_n2 & track_7_5_chanX_n5 & track_6_6_chanY_n13;
	track_6_5_chanX_n6_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_5_5_chanY_n6 & track_5_5_chanX_n6 & track_5_6_chanY_n5;
	track_6_5_chanX_n7_driver_mux_fanins  <= CLB_6_5_OUT_pin_2 & track_6_5_chanY_n4 & track_7_5_chanX_n7 & track_6_6_chanY_n11;
	track_6_5_chanX_n8_driver_mux_fanins  <= CLB_6_6_OUT_pin_0 & track_5_5_chanY_n4 & track_5_5_chanX_n8 & track_5_6_chanY_n7;
	track_6_5_chanX_n9_driver_mux_fanins  <= CLB_6_6_OUT_pin_0 & track_6_5_chanY_n6 & track_7_5_chanX_n9 & track_6_6_chanY_n9;
	track_6_5_chanY_n0_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_6_4_chanY_n0 & track_7_4_chanX_n3 & track_6_4_chanX_n0;
	track_6_5_chanY_n1_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_7_5_chanX_n13 & track_6_5_chanX_n2 & track_6_6_chanY_n1;
	track_6_5_chanY_n10_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_6_4_chanY_n10 & track_7_4_chanX_n13 & track_6_4_chanX_n6;
	track_6_5_chanY_n11_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_7_5_chanX_n3 & track_6_5_chanX_n12 & track_6_6_chanY_n11;
	track_6_5_chanY_n12_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_6_4_chanY_n12 & track_7_4_chanX_n15 & track_6_4_chanX_n4;
	track_6_5_chanY_n13_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_7_5_chanX_n1 & track_6_5_chanX_n14 & track_6_6_chanY_n13;
	track_6_5_chanY_n14_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_6_4_chanY_n14 & track_7_4_chanX_n1 & track_6_4_chanX_n2;
	track_6_5_chanY_n15_driver_mux_fanins <= CLB_7_5_OUT_pin_1 & track_7_5_chanX_n15 & track_6_5_chanX_n0 & track_6_6_chanY_n15;
	track_6_5_chanY_n2_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_6_4_chanY_n2 & track_7_4_chanX_n5 & track_6_4_chanX_n14;
	track_6_5_chanY_n3_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_7_5_chanX_n11 & track_6_5_chanX_n4 & track_6_6_chanY_n3;
	track_6_5_chanY_n4_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_6_4_chanY_n4 & track_7_4_chanX_n7 & track_6_4_chanX_n12;
	track_6_5_chanY_n5_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_7_5_chanX_n9 & track_6_5_chanX_n6 & track_6_6_chanY_n5;
	track_6_5_chanY_n6_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_6_4_chanY_n6 & track_7_4_chanX_n9 & track_6_4_chanX_n10;
	track_6_5_chanY_n7_driver_mux_fanins  <= CLB_6_5_OUT_pin_3 & track_7_5_chanX_n7 & track_6_5_chanX_n8 & track_6_6_chanY_n7;
	track_6_5_chanY_n8_driver_mux_fanins  <= CLB_7_5_OUT_pin_1 & track_6_4_chanY_n8 & track_7_4_chanX_n11 & track_6_4_chanX_n8;
	track_6_5_chanY_n9_driver_mux_fanins  <= CLB_7_5_OUT_pin_1 & track_7_5_chanX_n5 & track_6_5_chanX_n10 & track_6_6_chanY_n9;
	track_6_6_chanX_n0_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_5_6_chanY_n0 & track_5_6_chanX_n0;
	track_6_6_chanX_n1_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_6_6_chanY_n0 & track_7_6_chanX_n1;
	track_6_6_chanX_n10_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_5_6_chanY_n10 & track_5_6_chanX_n10;
	track_6_6_chanX_n11_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_6_6_chanY_n10 & track_7_6_chanX_n11;
	track_6_6_chanX_n12_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_5_6_chanY_n12 & track_5_6_chanX_n12;
	track_6_6_chanX_n13_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_6_6_chanY_n12 & track_7_6_chanX_n13;
	track_6_6_chanX_n14_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_5_6_chanY_n14 & track_5_6_chanX_n14;
	track_6_6_chanX_n15_driver_mux_fanins <= "0" & IO_6_7_OUT_pin_0 & track_6_6_chanY_n14 & track_7_6_chanX_n15;
	track_6_6_chanX_n2_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_5_6_chanY_n2 & track_5_6_chanX_n2;
	track_6_6_chanX_n3_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_6_6_chanY_n2 & track_7_6_chanX_n3;
	track_6_6_chanX_n4_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_5_6_chanY_n4 & track_5_6_chanX_n4;
	track_6_6_chanX_n5_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_6_6_chanY_n4 & track_7_6_chanX_n5;
	track_6_6_chanX_n6_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_5_6_chanY_n6 & track_5_6_chanX_n6;
	track_6_6_chanX_n7_driver_mux_fanins  <= IO_6_7_OUT_pin_1 & CLB_6_6_OUT_pin_2 & track_6_6_chanY_n6 & track_7_6_chanX_n7;
	track_6_6_chanX_n8_driver_mux_fanins  <= "0" & IO_6_7_OUT_pin_0 & track_5_6_chanY_n8 & track_5_6_chanX_n8;
	track_6_6_chanX_n9_driver_mux_fanins  <= "0" & IO_6_7_OUT_pin_0 & track_6_6_chanY_n8 & track_7_6_chanX_n9;
	track_6_6_chanY_n0_driver_mux_fanins  <= CLB_6_6_OUT_pin_3 & track_6_5_chanY_n0 & track_7_5_chanX_n3 & track_6_5_chanX_n0;
	track_6_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_6_6_OUT_pin_3 & track_7_6_chanX_n1 & track_6_6_chanX_n0;
	track_6_6_chanY_n10_driver_mux_fanins <= CLB_7_6_OUT_pin_1 & track_6_5_chanY_n10 & track_7_5_chanX_n13 & track_6_5_chanX_n6;
	track_6_6_chanY_n11_driver_mux_fanins <= "0" & CLB_7_6_OUT_pin_1 & track_7_6_chanX_n5 & track_6_6_chanX_n4;
	track_6_6_chanY_n12_driver_mux_fanins <= CLB_7_6_OUT_pin_1 & track_6_5_chanY_n12 & track_7_5_chanX_n15 & track_6_5_chanX_n4;
	track_6_6_chanY_n13_driver_mux_fanins <= "0" & CLB_7_6_OUT_pin_1 & track_7_6_chanX_n7 & track_6_6_chanX_n6;
	track_6_6_chanY_n14_driver_mux_fanins <= CLB_7_6_OUT_pin_1 & track_6_5_chanY_n14 & track_7_5_chanX_n1 & track_6_5_chanX_n2;
	track_6_6_chanY_n15_driver_mux_fanins <= "0" & CLB_7_6_OUT_pin_1 & track_7_6_chanX_n15 & track_6_6_chanX_n14;
	track_6_6_chanY_n2_driver_mux_fanins  <= CLB_6_6_OUT_pin_3 & track_6_5_chanY_n2 & track_7_5_chanX_n5 & track_6_5_chanX_n14;
	track_6_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_6_6_OUT_pin_3 & track_7_6_chanX_n9 & track_6_6_chanX_n8;
	track_6_6_chanY_n4_driver_mux_fanins  <= CLB_6_6_OUT_pin_3 & track_6_5_chanY_n4 & track_7_5_chanX_n7 & track_6_5_chanX_n12;
	track_6_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_6_6_OUT_pin_3 & track_7_6_chanX_n11 & track_6_6_chanX_n10;
	track_6_6_chanY_n6_driver_mux_fanins  <= CLB_6_6_OUT_pin_3 & track_6_5_chanY_n6 & track_7_5_chanX_n9 & track_6_5_chanX_n10;
	track_6_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_6_6_OUT_pin_3 & track_7_6_chanX_n13 & track_6_6_chanX_n12;
	track_6_6_chanY_n8_driver_mux_fanins  <= CLB_7_6_OUT_pin_1 & track_6_5_chanY_n8 & track_7_5_chanX_n11 & track_6_5_chanX_n8;
	track_6_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_7_6_OUT_pin_1 & track_7_6_chanX_n3 & track_6_6_chanX_n2;
	track_7_0_chanX_n0_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_6_0_chanX_n0 & track_6_1_chanY_n1;
	track_7_0_chanX_n1_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_8_0_chanX_n1 & track_7_1_chanY_n1;
	track_7_0_chanX_n10_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_6_0_chanX_n10 & track_6_1_chanY_n11;
	track_7_0_chanX_n11_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_8_0_chanX_n11 & track_7_1_chanY_n11;
	track_7_0_chanX_n12_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_6_0_chanX_n12 & track_6_1_chanY_n13;
	track_7_0_chanX_n13_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_8_0_chanX_n13 & track_7_1_chanY_n13;
	track_7_0_chanX_n14_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_6_0_chanX_n14 & track_6_1_chanY_n15;
	track_7_0_chanX_n15_driver_mux_fanins <= "0" & IO_7_0_OUT_pin_1 & track_8_0_chanX_n15 & track_7_1_chanY_n15;
	track_7_0_chanX_n2_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_6_0_chanX_n2 & track_6_1_chanY_n3;
	track_7_0_chanX_n3_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_8_0_chanX_n3 & track_7_1_chanY_n3;
	track_7_0_chanX_n4_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_6_0_chanX_n4 & track_6_1_chanY_n5;
	track_7_0_chanX_n5_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_8_0_chanX_n5 & track_7_1_chanY_n5;
	track_7_0_chanX_n6_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_6_0_chanX_n6 & track_6_1_chanY_n7;
	track_7_0_chanX_n7_driver_mux_fanins  <= IO_7_0_OUT_pin_0 & CLB_7_1_OUT_pin_0 & track_8_0_chanX_n7 & track_7_1_chanY_n7;
	track_7_0_chanX_n8_driver_mux_fanins  <= "0" & IO_7_0_OUT_pin_1 & track_6_0_chanX_n8 & track_6_1_chanY_n9;
	track_7_0_chanX_n9_driver_mux_fanins  <= "0" & IO_7_0_OUT_pin_1 & track_8_0_chanX_n9 & track_7_1_chanY_n9;
	track_7_1_chanX_n0_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_6_1_chanY_n12 & track_6_1_chanX_n0 & track_6_2_chanY_n15;
	track_7_1_chanX_n1_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_7_1_chanY_n14 & track_8_1_chanX_n1 & track_7_2_chanY_n1;
	track_7_1_chanX_n10_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_6_1_chanY_n2 & track_6_1_chanX_n10 & track_6_2_chanY_n9;
	track_7_1_chanX_n11_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_7_1_chanY_n8 & track_8_1_chanX_n11 & track_7_2_chanY_n7;
	track_7_1_chanX_n12_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_6_1_chanY_n0 & track_6_1_chanX_n12 & track_6_2_chanY_n11;
	track_7_1_chanX_n13_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_7_1_chanY_n10 & track_8_1_chanX_n13 & track_7_2_chanY_n5;
	track_7_1_chanX_n14_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_6_1_chanY_n14 & track_6_1_chanX_n14 & track_6_2_chanY_n13;
	track_7_1_chanX_n15_driver_mux_fanins <= CLB_7_2_OUT_pin_0 & track_7_1_chanY_n12 & track_8_1_chanX_n15 & track_7_2_chanY_n3;
	track_7_1_chanX_n2_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_6_1_chanY_n10 & track_6_1_chanX_n2 & track_6_2_chanY_n1;
	track_7_1_chanX_n3_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_7_1_chanY_n0 & track_8_1_chanX_n3 & track_7_2_chanY_n15;
	track_7_1_chanX_n4_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_6_1_chanY_n8 & track_6_1_chanX_n4 & track_6_2_chanY_n3;
	track_7_1_chanX_n5_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_7_1_chanY_n2 & track_8_1_chanX_n5 & track_7_2_chanY_n13;
	track_7_1_chanX_n6_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_6_1_chanY_n6 & track_6_1_chanX_n6 & track_6_2_chanY_n5;
	track_7_1_chanX_n7_driver_mux_fanins  <= CLB_7_1_OUT_pin_2 & track_7_1_chanY_n4 & track_8_1_chanX_n7 & track_7_2_chanY_n11;
	track_7_1_chanX_n8_driver_mux_fanins  <= CLB_7_2_OUT_pin_0 & track_6_1_chanY_n4 & track_6_1_chanX_n8 & track_6_2_chanY_n7;
	track_7_1_chanX_n9_driver_mux_fanins  <= CLB_7_2_OUT_pin_0 & track_7_1_chanY_n6 & track_8_1_chanX_n9 & track_7_2_chanY_n9;
	track_7_1_chanY_n0_driver_mux_fanins  <= "0" & CLB_7_1_OUT_pin_3 & track_8_0_chanX_n7 & track_7_0_chanX_n6;
	track_7_1_chanY_n1_driver_mux_fanins  <= CLB_7_1_OUT_pin_3 & track_8_1_chanX_n13 & track_7_1_chanX_n2 & track_7_2_chanY_n1;
	track_7_1_chanY_n10_driver_mux_fanins <= "0" & CLB_8_1_OUT_pin_1 & track_8_0_chanX_n11 & track_7_0_chanX_n10;
	track_7_1_chanY_n11_driver_mux_fanins <= CLB_8_1_OUT_pin_1 & track_8_1_chanX_n3 & track_7_1_chanX_n12 & track_7_2_chanY_n11;
	track_7_1_chanY_n12_driver_mux_fanins <= "0" & CLB_8_1_OUT_pin_1 & track_8_0_chanX_n13 & track_7_0_chanX_n12;
	track_7_1_chanY_n13_driver_mux_fanins <= CLB_8_1_OUT_pin_1 & track_8_1_chanX_n1 & track_7_1_chanX_n14 & track_7_2_chanY_n13;
	track_7_1_chanY_n14_driver_mux_fanins <= "0" & CLB_8_1_OUT_pin_1 & track_8_0_chanX_n15 & track_7_0_chanX_n14;
	track_7_1_chanY_n15_driver_mux_fanins <= CLB_8_1_OUT_pin_1 & track_8_1_chanX_n15 & track_7_1_chanX_n0 & track_7_2_chanY_n15;
	track_7_1_chanY_n2_driver_mux_fanins  <= "0" & CLB_7_1_OUT_pin_3 & track_8_0_chanX_n9 & track_7_0_chanX_n8;
	track_7_1_chanY_n3_driver_mux_fanins  <= CLB_7_1_OUT_pin_3 & track_8_1_chanX_n11 & track_7_1_chanX_n4 & track_7_2_chanY_n3;
	track_7_1_chanY_n4_driver_mux_fanins  <= "0" & CLB_7_1_OUT_pin_3 & track_8_0_chanX_n1 & track_7_0_chanX_n0;
	track_7_1_chanY_n5_driver_mux_fanins  <= CLB_7_1_OUT_pin_3 & track_8_1_chanX_n9 & track_7_1_chanX_n6 & track_7_2_chanY_n5;
	track_7_1_chanY_n6_driver_mux_fanins  <= "0" & CLB_7_1_OUT_pin_3 & track_8_0_chanX_n3 & track_7_0_chanX_n2;
	track_7_1_chanY_n7_driver_mux_fanins  <= CLB_7_1_OUT_pin_3 & track_8_1_chanX_n7 & track_7_1_chanX_n8 & track_7_2_chanY_n7;
	track_7_1_chanY_n8_driver_mux_fanins  <= "0" & CLB_8_1_OUT_pin_1 & track_8_0_chanX_n5 & track_7_0_chanX_n4;
	track_7_1_chanY_n9_driver_mux_fanins  <= CLB_8_1_OUT_pin_1 & track_8_1_chanX_n5 & track_7_1_chanX_n10 & track_7_2_chanY_n9;
	track_7_2_chanX_n0_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_6_2_chanY_n12 & track_6_2_chanX_n0 & track_6_3_chanY_n15;
	track_7_2_chanX_n1_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_7_2_chanY_n14 & track_8_2_chanX_n1 & track_7_3_chanY_n1;
	track_7_2_chanX_n10_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_6_2_chanY_n2 & track_6_2_chanX_n10 & track_6_3_chanY_n9;
	track_7_2_chanX_n11_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_7_2_chanY_n8 & track_8_2_chanX_n11 & track_7_3_chanY_n7;
	track_7_2_chanX_n12_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_6_2_chanY_n0 & track_6_2_chanX_n12 & track_6_3_chanY_n11;
	track_7_2_chanX_n13_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_7_2_chanY_n10 & track_8_2_chanX_n13 & track_7_3_chanY_n5;
	track_7_2_chanX_n14_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_6_2_chanY_n14 & track_6_2_chanX_n14 & track_6_3_chanY_n13;
	track_7_2_chanX_n15_driver_mux_fanins <= CLB_7_3_OUT_pin_0 & track_7_2_chanY_n12 & track_8_2_chanX_n15 & track_7_3_chanY_n3;
	track_7_2_chanX_n2_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_6_2_chanY_n10 & track_6_2_chanX_n2 & track_6_3_chanY_n1;
	track_7_2_chanX_n3_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_7_2_chanY_n0 & track_8_2_chanX_n3 & track_7_3_chanY_n15;
	track_7_2_chanX_n4_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_6_2_chanY_n8 & track_6_2_chanX_n4 & track_6_3_chanY_n3;
	track_7_2_chanX_n5_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_7_2_chanY_n2 & track_8_2_chanX_n5 & track_7_3_chanY_n13;
	track_7_2_chanX_n6_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_6_2_chanY_n6 & track_6_2_chanX_n6 & track_6_3_chanY_n5;
	track_7_2_chanX_n7_driver_mux_fanins  <= CLB_7_2_OUT_pin_2 & track_7_2_chanY_n4 & track_8_2_chanX_n7 & track_7_3_chanY_n11;
	track_7_2_chanX_n8_driver_mux_fanins  <= CLB_7_3_OUT_pin_0 & track_6_2_chanY_n4 & track_6_2_chanX_n8 & track_6_3_chanY_n7;
	track_7_2_chanX_n9_driver_mux_fanins  <= CLB_7_3_OUT_pin_0 & track_7_2_chanY_n6 & track_8_2_chanX_n9 & track_7_3_chanY_n9;
	track_7_2_chanY_n0_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_7_1_chanY_n0 & track_8_1_chanX_n3 & track_7_1_chanX_n0;
	track_7_2_chanY_n1_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_8_2_chanX_n13 & track_7_2_chanX_n2 & track_7_3_chanY_n1;
	track_7_2_chanY_n10_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_7_1_chanY_n10 & track_8_1_chanX_n13 & track_7_1_chanX_n6;
	track_7_2_chanY_n11_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_8_2_chanX_n3 & track_7_2_chanX_n12 & track_7_3_chanY_n11;
	track_7_2_chanY_n12_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_7_1_chanY_n12 & track_8_1_chanX_n15 & track_7_1_chanX_n4;
	track_7_2_chanY_n13_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_8_2_chanX_n1 & track_7_2_chanX_n14 & track_7_3_chanY_n13;
	track_7_2_chanY_n14_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_7_1_chanY_n14 & track_8_1_chanX_n1 & track_7_1_chanX_n2;
	track_7_2_chanY_n15_driver_mux_fanins <= CLB_8_2_OUT_pin_1 & track_8_2_chanX_n15 & track_7_2_chanX_n0 & track_7_3_chanY_n15;
	track_7_2_chanY_n2_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_7_1_chanY_n2 & track_8_1_chanX_n5 & track_7_1_chanX_n14;
	track_7_2_chanY_n3_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_8_2_chanX_n11 & track_7_2_chanX_n4 & track_7_3_chanY_n3;
	track_7_2_chanY_n4_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_7_1_chanY_n4 & track_8_1_chanX_n7 & track_7_1_chanX_n12;
	track_7_2_chanY_n5_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_8_2_chanX_n9 & track_7_2_chanX_n6 & track_7_3_chanY_n5;
	track_7_2_chanY_n6_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_7_1_chanY_n6 & track_8_1_chanX_n9 & track_7_1_chanX_n10;
	track_7_2_chanY_n7_driver_mux_fanins  <= CLB_7_2_OUT_pin_3 & track_8_2_chanX_n7 & track_7_2_chanX_n8 & track_7_3_chanY_n7;
	track_7_2_chanY_n8_driver_mux_fanins  <= CLB_8_2_OUT_pin_1 & track_7_1_chanY_n8 & track_8_1_chanX_n11 & track_7_1_chanX_n8;
	track_7_2_chanY_n9_driver_mux_fanins  <= CLB_8_2_OUT_pin_1 & track_8_2_chanX_n5 & track_7_2_chanX_n10 & track_7_3_chanY_n9;
	track_7_3_chanX_n0_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_6_3_chanY_n12 & track_6_3_chanX_n0 & track_6_4_chanY_n15;
	track_7_3_chanX_n1_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_7_3_chanY_n14 & track_8_3_chanX_n1 & track_7_4_chanY_n1;
	track_7_3_chanX_n10_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_6_3_chanY_n2 & track_6_3_chanX_n10 & track_6_4_chanY_n9;
	track_7_3_chanX_n11_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_7_3_chanY_n8 & track_8_3_chanX_n11 & track_7_4_chanY_n7;
	track_7_3_chanX_n12_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_6_3_chanY_n0 & track_6_3_chanX_n12 & track_6_4_chanY_n11;
	track_7_3_chanX_n13_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_7_3_chanY_n10 & track_8_3_chanX_n13 & track_7_4_chanY_n5;
	track_7_3_chanX_n14_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_6_3_chanY_n14 & track_6_3_chanX_n14 & track_6_4_chanY_n13;
	track_7_3_chanX_n15_driver_mux_fanins <= CLB_7_4_OUT_pin_0 & track_7_3_chanY_n12 & track_8_3_chanX_n15 & track_7_4_chanY_n3;
	track_7_3_chanX_n2_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_6_3_chanY_n10 & track_6_3_chanX_n2 & track_6_4_chanY_n1;
	track_7_3_chanX_n3_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_7_3_chanY_n0 & track_8_3_chanX_n3 & track_7_4_chanY_n15;
	track_7_3_chanX_n4_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_6_3_chanY_n8 & track_6_3_chanX_n4 & track_6_4_chanY_n3;
	track_7_3_chanX_n5_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_7_3_chanY_n2 & track_8_3_chanX_n5 & track_7_4_chanY_n13;
	track_7_3_chanX_n6_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_6_3_chanY_n6 & track_6_3_chanX_n6 & track_6_4_chanY_n5;
	track_7_3_chanX_n7_driver_mux_fanins  <= CLB_7_3_OUT_pin_2 & track_7_3_chanY_n4 & track_8_3_chanX_n7 & track_7_4_chanY_n11;
	track_7_3_chanX_n8_driver_mux_fanins  <= CLB_7_4_OUT_pin_0 & track_6_3_chanY_n4 & track_6_3_chanX_n8 & track_6_4_chanY_n7;
	track_7_3_chanX_n9_driver_mux_fanins  <= CLB_7_4_OUT_pin_0 & track_7_3_chanY_n6 & track_8_3_chanX_n9 & track_7_4_chanY_n9;
	track_7_3_chanY_n0_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_7_2_chanY_n0 & track_8_2_chanX_n3 & track_7_2_chanX_n0;
	track_7_3_chanY_n1_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_8_3_chanX_n13 & track_7_3_chanX_n2 & track_7_4_chanY_n1;
	track_7_3_chanY_n10_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_7_2_chanY_n10 & track_8_2_chanX_n13 & track_7_2_chanX_n6;
	track_7_3_chanY_n11_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_8_3_chanX_n3 & track_7_3_chanX_n12 & track_7_4_chanY_n11;
	track_7_3_chanY_n12_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_7_2_chanY_n12 & track_8_2_chanX_n15 & track_7_2_chanX_n4;
	track_7_3_chanY_n13_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_8_3_chanX_n1 & track_7_3_chanX_n14 & track_7_4_chanY_n13;
	track_7_3_chanY_n14_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_7_2_chanY_n14 & track_8_2_chanX_n1 & track_7_2_chanX_n2;
	track_7_3_chanY_n15_driver_mux_fanins <= CLB_8_3_OUT_pin_1 & track_8_3_chanX_n15 & track_7_3_chanX_n0 & track_7_4_chanY_n15;
	track_7_3_chanY_n2_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_7_2_chanY_n2 & track_8_2_chanX_n5 & track_7_2_chanX_n14;
	track_7_3_chanY_n3_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_8_3_chanX_n11 & track_7_3_chanX_n4 & track_7_4_chanY_n3;
	track_7_3_chanY_n4_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_7_2_chanY_n4 & track_8_2_chanX_n7 & track_7_2_chanX_n12;
	track_7_3_chanY_n5_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_8_3_chanX_n9 & track_7_3_chanX_n6 & track_7_4_chanY_n5;
	track_7_3_chanY_n6_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_7_2_chanY_n6 & track_8_2_chanX_n9 & track_7_2_chanX_n10;
	track_7_3_chanY_n7_driver_mux_fanins  <= CLB_7_3_OUT_pin_3 & track_8_3_chanX_n7 & track_7_3_chanX_n8 & track_7_4_chanY_n7;
	track_7_3_chanY_n8_driver_mux_fanins  <= CLB_8_3_OUT_pin_1 & track_7_2_chanY_n8 & track_8_2_chanX_n11 & track_7_2_chanX_n8;
	track_7_3_chanY_n9_driver_mux_fanins  <= CLB_8_3_OUT_pin_1 & track_8_3_chanX_n5 & track_7_3_chanX_n10 & track_7_4_chanY_n9;
	track_7_4_chanX_n0_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_6_4_chanY_n12 & track_6_4_chanX_n0 & track_6_5_chanY_n15;
	track_7_4_chanX_n1_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_7_4_chanY_n14 & track_8_4_chanX_n1 & track_7_5_chanY_n1;
	track_7_4_chanX_n10_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_6_4_chanY_n2 & track_6_4_chanX_n10 & track_6_5_chanY_n9;
	track_7_4_chanX_n11_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_7_4_chanY_n8 & track_8_4_chanX_n11 & track_7_5_chanY_n7;
	track_7_4_chanX_n12_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_6_4_chanY_n0 & track_6_4_chanX_n12 & track_6_5_chanY_n11;
	track_7_4_chanX_n13_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_7_4_chanY_n10 & track_8_4_chanX_n13 & track_7_5_chanY_n5;
	track_7_4_chanX_n14_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_6_4_chanY_n14 & track_6_4_chanX_n14 & track_6_5_chanY_n13;
	track_7_4_chanX_n15_driver_mux_fanins <= CLB_7_5_OUT_pin_0 & track_7_4_chanY_n12 & track_8_4_chanX_n15 & track_7_5_chanY_n3;
	track_7_4_chanX_n2_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_6_4_chanY_n10 & track_6_4_chanX_n2 & track_6_5_chanY_n1;
	track_7_4_chanX_n3_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_7_4_chanY_n0 & track_8_4_chanX_n3 & track_7_5_chanY_n15;
	track_7_4_chanX_n4_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_6_4_chanY_n8 & track_6_4_chanX_n4 & track_6_5_chanY_n3;
	track_7_4_chanX_n5_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_7_4_chanY_n2 & track_8_4_chanX_n5 & track_7_5_chanY_n13;
	track_7_4_chanX_n6_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_6_4_chanY_n6 & track_6_4_chanX_n6 & track_6_5_chanY_n5;
	track_7_4_chanX_n7_driver_mux_fanins  <= CLB_7_4_OUT_pin_2 & track_7_4_chanY_n4 & track_8_4_chanX_n7 & track_7_5_chanY_n11;
	track_7_4_chanX_n8_driver_mux_fanins  <= CLB_7_5_OUT_pin_0 & track_6_4_chanY_n4 & track_6_4_chanX_n8 & track_6_5_chanY_n7;
	track_7_4_chanX_n9_driver_mux_fanins  <= CLB_7_5_OUT_pin_0 & track_7_4_chanY_n6 & track_8_4_chanX_n9 & track_7_5_chanY_n9;
	track_7_4_chanY_n0_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_7_3_chanY_n0 & track_8_3_chanX_n3 & track_7_3_chanX_n0;
	track_7_4_chanY_n1_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_8_4_chanX_n13 & track_7_4_chanX_n2 & track_7_5_chanY_n1;
	track_7_4_chanY_n10_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_7_3_chanY_n10 & track_8_3_chanX_n13 & track_7_3_chanX_n6;
	track_7_4_chanY_n11_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_8_4_chanX_n3 & track_7_4_chanX_n12 & track_7_5_chanY_n11;
	track_7_4_chanY_n12_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_7_3_chanY_n12 & track_8_3_chanX_n15 & track_7_3_chanX_n4;
	track_7_4_chanY_n13_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_8_4_chanX_n1 & track_7_4_chanX_n14 & track_7_5_chanY_n13;
	track_7_4_chanY_n14_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_7_3_chanY_n14 & track_8_3_chanX_n1 & track_7_3_chanX_n2;
	track_7_4_chanY_n15_driver_mux_fanins <= CLB_8_4_OUT_pin_1 & track_8_4_chanX_n15 & track_7_4_chanX_n0 & track_7_5_chanY_n15;
	track_7_4_chanY_n2_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_7_3_chanY_n2 & track_8_3_chanX_n5 & track_7_3_chanX_n14;
	track_7_4_chanY_n3_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_8_4_chanX_n11 & track_7_4_chanX_n4 & track_7_5_chanY_n3;
	track_7_4_chanY_n4_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_7_3_chanY_n4 & track_8_3_chanX_n7 & track_7_3_chanX_n12;
	track_7_4_chanY_n5_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_8_4_chanX_n9 & track_7_4_chanX_n6 & track_7_5_chanY_n5;
	track_7_4_chanY_n6_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_7_3_chanY_n6 & track_8_3_chanX_n9 & track_7_3_chanX_n10;
	track_7_4_chanY_n7_driver_mux_fanins  <= CLB_7_4_OUT_pin_3 & track_8_4_chanX_n7 & track_7_4_chanX_n8 & track_7_5_chanY_n7;
	track_7_4_chanY_n8_driver_mux_fanins  <= CLB_8_4_OUT_pin_1 & track_7_3_chanY_n8 & track_8_3_chanX_n11 & track_7_3_chanX_n8;
	track_7_4_chanY_n9_driver_mux_fanins  <= CLB_8_4_OUT_pin_1 & track_8_4_chanX_n5 & track_7_4_chanX_n10 & track_7_5_chanY_n9;
	track_7_5_chanX_n0_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_6_5_chanY_n12 & track_6_5_chanX_n0 & track_6_6_chanY_n15;
	track_7_5_chanX_n1_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_7_5_chanY_n14 & track_8_5_chanX_n1 & track_7_6_chanY_n1;
	track_7_5_chanX_n10_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_6_5_chanY_n2 & track_6_5_chanX_n10 & track_6_6_chanY_n9;
	track_7_5_chanX_n11_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_7_5_chanY_n8 & track_8_5_chanX_n11 & track_7_6_chanY_n7;
	track_7_5_chanX_n12_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_6_5_chanY_n0 & track_6_5_chanX_n12 & track_6_6_chanY_n11;
	track_7_5_chanX_n13_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_7_5_chanY_n10 & track_8_5_chanX_n13 & track_7_6_chanY_n5;
	track_7_5_chanX_n14_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_6_5_chanY_n14 & track_6_5_chanX_n14 & track_6_6_chanY_n13;
	track_7_5_chanX_n15_driver_mux_fanins <= CLB_7_6_OUT_pin_0 & track_7_5_chanY_n12 & track_8_5_chanX_n15 & track_7_6_chanY_n3;
	track_7_5_chanX_n2_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_6_5_chanY_n10 & track_6_5_chanX_n2 & track_6_6_chanY_n1;
	track_7_5_chanX_n3_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_7_5_chanY_n0 & track_8_5_chanX_n3 & track_7_6_chanY_n15;
	track_7_5_chanX_n4_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_6_5_chanY_n8 & track_6_5_chanX_n4 & track_6_6_chanY_n3;
	track_7_5_chanX_n5_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_7_5_chanY_n2 & track_8_5_chanX_n5 & track_7_6_chanY_n13;
	track_7_5_chanX_n6_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_6_5_chanY_n6 & track_6_5_chanX_n6 & track_6_6_chanY_n5;
	track_7_5_chanX_n7_driver_mux_fanins  <= CLB_7_5_OUT_pin_2 & track_7_5_chanY_n4 & track_8_5_chanX_n7 & track_7_6_chanY_n11;
	track_7_5_chanX_n8_driver_mux_fanins  <= CLB_7_6_OUT_pin_0 & track_6_5_chanY_n4 & track_6_5_chanX_n8 & track_6_6_chanY_n7;
	track_7_5_chanX_n9_driver_mux_fanins  <= CLB_7_6_OUT_pin_0 & track_7_5_chanY_n6 & track_8_5_chanX_n9 & track_7_6_chanY_n9;
	track_7_5_chanY_n0_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_7_4_chanY_n0 & track_8_4_chanX_n3 & track_7_4_chanX_n0;
	track_7_5_chanY_n1_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_8_5_chanX_n13 & track_7_5_chanX_n2 & track_7_6_chanY_n1;
	track_7_5_chanY_n10_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_7_4_chanY_n10 & track_8_4_chanX_n13 & track_7_4_chanX_n6;
	track_7_5_chanY_n11_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_8_5_chanX_n3 & track_7_5_chanX_n12 & track_7_6_chanY_n11;
	track_7_5_chanY_n12_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_7_4_chanY_n12 & track_8_4_chanX_n15 & track_7_4_chanX_n4;
	track_7_5_chanY_n13_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_8_5_chanX_n1 & track_7_5_chanX_n14 & track_7_6_chanY_n13;
	track_7_5_chanY_n14_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_7_4_chanY_n14 & track_8_4_chanX_n1 & track_7_4_chanX_n2;
	track_7_5_chanY_n15_driver_mux_fanins <= CLB_8_5_OUT_pin_1 & track_8_5_chanX_n15 & track_7_5_chanX_n0 & track_7_6_chanY_n15;
	track_7_5_chanY_n2_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_7_4_chanY_n2 & track_8_4_chanX_n5 & track_7_4_chanX_n14;
	track_7_5_chanY_n3_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_8_5_chanX_n11 & track_7_5_chanX_n4 & track_7_6_chanY_n3;
	track_7_5_chanY_n4_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_7_4_chanY_n4 & track_8_4_chanX_n7 & track_7_4_chanX_n12;
	track_7_5_chanY_n5_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_8_5_chanX_n9 & track_7_5_chanX_n6 & track_7_6_chanY_n5;
	track_7_5_chanY_n6_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_7_4_chanY_n6 & track_8_4_chanX_n9 & track_7_4_chanX_n10;
	track_7_5_chanY_n7_driver_mux_fanins  <= CLB_7_5_OUT_pin_3 & track_8_5_chanX_n7 & track_7_5_chanX_n8 & track_7_6_chanY_n7;
	track_7_5_chanY_n8_driver_mux_fanins  <= CLB_8_5_OUT_pin_1 & track_7_4_chanY_n8 & track_8_4_chanX_n11 & track_7_4_chanX_n8;
	track_7_5_chanY_n9_driver_mux_fanins  <= CLB_8_5_OUT_pin_1 & track_8_5_chanX_n5 & track_7_5_chanX_n10 & track_7_6_chanY_n9;
	track_7_6_chanX_n0_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_6_6_chanY_n0 & track_6_6_chanX_n0;
	track_7_6_chanX_n1_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_7_6_chanY_n0 & track_8_6_chanX_n1;
	track_7_6_chanX_n10_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_6_6_chanY_n10 & track_6_6_chanX_n10;
	track_7_6_chanX_n11_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_7_6_chanY_n10 & track_8_6_chanX_n11;
	track_7_6_chanX_n12_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_6_6_chanY_n12 & track_6_6_chanX_n12;
	track_7_6_chanX_n13_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_7_6_chanY_n12 & track_8_6_chanX_n13;
	track_7_6_chanX_n14_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_6_6_chanY_n14 & track_6_6_chanX_n14;
	track_7_6_chanX_n15_driver_mux_fanins <= "0" & IO_7_7_OUT_pin_0 & track_7_6_chanY_n14 & track_8_6_chanX_n15;
	track_7_6_chanX_n2_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_6_6_chanY_n2 & track_6_6_chanX_n2;
	track_7_6_chanX_n3_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_7_6_chanY_n2 & track_8_6_chanX_n3;
	track_7_6_chanX_n4_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_6_6_chanY_n4 & track_6_6_chanX_n4;
	track_7_6_chanX_n5_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_7_6_chanY_n4 & track_8_6_chanX_n5;
	track_7_6_chanX_n6_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_6_6_chanY_n6 & track_6_6_chanX_n6;
	track_7_6_chanX_n7_driver_mux_fanins  <= IO_7_7_OUT_pin_1 & CLB_7_6_OUT_pin_2 & track_7_6_chanY_n6 & track_8_6_chanX_n7;
	track_7_6_chanX_n8_driver_mux_fanins  <= "0" & IO_7_7_OUT_pin_0 & track_6_6_chanY_n8 & track_6_6_chanX_n8;
	track_7_6_chanX_n9_driver_mux_fanins  <= "0" & IO_7_7_OUT_pin_0 & track_7_6_chanY_n8 & track_8_6_chanX_n9;
	track_7_6_chanY_n0_driver_mux_fanins  <= CLB_7_6_OUT_pin_3 & track_7_5_chanY_n0 & track_8_5_chanX_n3 & track_7_5_chanX_n0;
	track_7_6_chanY_n1_driver_mux_fanins  <= "0" & CLB_7_6_OUT_pin_3 & track_8_6_chanX_n1 & track_7_6_chanX_n0;
	track_7_6_chanY_n10_driver_mux_fanins <= CLB_8_6_OUT_pin_1 & track_7_5_chanY_n10 & track_8_5_chanX_n13 & track_7_5_chanX_n6;
	track_7_6_chanY_n11_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_1 & track_8_6_chanX_n5 & track_7_6_chanX_n4;
	track_7_6_chanY_n12_driver_mux_fanins <= CLB_8_6_OUT_pin_1 & track_7_5_chanY_n12 & track_8_5_chanX_n15 & track_7_5_chanX_n4;
	track_7_6_chanY_n13_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_1 & track_8_6_chanX_n7 & track_7_6_chanX_n6;
	track_7_6_chanY_n14_driver_mux_fanins <= CLB_8_6_OUT_pin_1 & track_7_5_chanY_n14 & track_8_5_chanX_n1 & track_7_5_chanX_n2;
	track_7_6_chanY_n15_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_1 & track_8_6_chanX_n15 & track_7_6_chanX_n14;
	track_7_6_chanY_n2_driver_mux_fanins  <= CLB_7_6_OUT_pin_3 & track_7_5_chanY_n2 & track_8_5_chanX_n5 & track_7_5_chanX_n14;
	track_7_6_chanY_n3_driver_mux_fanins  <= "0" & CLB_7_6_OUT_pin_3 & track_8_6_chanX_n9 & track_7_6_chanX_n8;
	track_7_6_chanY_n4_driver_mux_fanins  <= CLB_7_6_OUT_pin_3 & track_7_5_chanY_n4 & track_8_5_chanX_n7 & track_7_5_chanX_n12;
	track_7_6_chanY_n5_driver_mux_fanins  <= "0" & CLB_7_6_OUT_pin_3 & track_8_6_chanX_n11 & track_7_6_chanX_n10;
	track_7_6_chanY_n6_driver_mux_fanins  <= CLB_7_6_OUT_pin_3 & track_7_5_chanY_n6 & track_8_5_chanX_n9 & track_7_5_chanX_n10;
	track_7_6_chanY_n7_driver_mux_fanins  <= "0" & CLB_7_6_OUT_pin_3 & track_8_6_chanX_n13 & track_7_6_chanX_n12;
	track_7_6_chanY_n8_driver_mux_fanins  <= CLB_8_6_OUT_pin_1 & track_7_5_chanY_n8 & track_8_5_chanX_n11 & track_7_5_chanX_n8;
	track_7_6_chanY_n9_driver_mux_fanins  <= "0" & CLB_8_6_OUT_pin_1 & track_8_6_chanX_n3 & track_7_6_chanX_n2;
	track_8_0_chanX_n0_driver_mux_fanins  <= IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_7_0_chanX_n0 & track_7_1_chanY_n1;
	track_8_0_chanX_n1_driver_mux_fanins  <= "0" & IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_8_1_chanY_n1;
	track_8_0_chanX_n10_driver_mux_fanins <= "0" & IO_8_0_OUT_pin_1 & track_7_0_chanX_n10 & track_7_1_chanY_n11;
	track_8_0_chanX_n11_driver_mux_fanins <= IO_8_0_OUT_pin_1 & track_8_1_chanY_n7;
	track_8_0_chanX_n12_driver_mux_fanins <= "0" & IO_8_0_OUT_pin_1 & track_7_0_chanX_n12 & track_7_1_chanY_n13;
	track_8_0_chanX_n13_driver_mux_fanins <= IO_8_0_OUT_pin_1 & track_8_1_chanY_n5;
	track_8_0_chanX_n14_driver_mux_fanins <= "0" & IO_8_0_OUT_pin_1 & track_7_0_chanX_n14 & track_7_1_chanY_n15;
	track_8_0_chanX_n15_driver_mux_fanins <= IO_8_0_OUT_pin_1 & track_8_1_chanY_n3;
	track_8_0_chanX_n2_driver_mux_fanins  <= IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_7_0_chanX_n2 & track_7_1_chanY_n3;
	track_8_0_chanX_n3_driver_mux_fanins  <= "0" & IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_8_1_chanY_n15;
	track_8_0_chanX_n4_driver_mux_fanins  <= IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_7_0_chanX_n4 & track_7_1_chanY_n5;
	track_8_0_chanX_n5_driver_mux_fanins  <= "0" & IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_8_1_chanY_n13;
	track_8_0_chanX_n6_driver_mux_fanins  <= IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_7_0_chanX_n6 & track_7_1_chanY_n7;
	track_8_0_chanX_n7_driver_mux_fanins  <= "0" & IO_8_0_OUT_pin_0 & CLB_8_1_OUT_pin_0 & track_8_1_chanY_n11;
	track_8_0_chanX_n8_driver_mux_fanins  <= "0" & IO_8_0_OUT_pin_1 & track_7_0_chanX_n8 & track_7_1_chanY_n9;
	track_8_0_chanX_n9_driver_mux_fanins  <= IO_8_0_OUT_pin_1 & track_8_1_chanY_n9;
	track_8_1_chanX_n0_driver_mux_fanins  <= CLB_8_1_OUT_pin_2 & track_7_1_chanY_n12 & track_7_1_chanX_n0 & track_7_2_chanY_n15;
	track_8_1_chanX_n1_driver_mux_fanins  <= "0" & CLB_8_1_OUT_pin_2 & track_8_1_chanY_n0 & track_8_2_chanY_n1;
	track_8_1_chanX_n10_driver_mux_fanins <= CLB_8_2_OUT_pin_0 & track_7_1_chanY_n2 & track_7_1_chanX_n10 & track_7_2_chanY_n9;
	track_8_1_chanX_n11_driver_mux_fanins <= "0" & CLB_8_2_OUT_pin_0 & track_8_1_chanY_n4 & track_8_2_chanY_n5;
	track_8_1_chanX_n12_driver_mux_fanins <= CLB_8_2_OUT_pin_0 & track_7_1_chanY_n0 & track_7_1_chanX_n12 & track_7_2_chanY_n11;
	track_8_1_chanX_n13_driver_mux_fanins <= "0" & CLB_8_2_OUT_pin_0 & track_8_1_chanY_n6 & track_8_2_chanY_n7;
	track_8_1_chanX_n14_driver_mux_fanins <= CLB_8_2_OUT_pin_0 & track_7_1_chanY_n14 & track_7_1_chanX_n14 & track_7_2_chanY_n13;
	track_8_1_chanX_n15_driver_mux_fanins <= "0" & CLB_8_2_OUT_pin_0 & track_8_1_chanY_n14 & track_8_2_chanY_n15;
	track_8_1_chanX_n2_driver_mux_fanins  <= CLB_8_1_OUT_pin_2 & track_7_1_chanY_n10 & track_7_1_chanX_n2 & track_7_2_chanY_n1;
	track_8_1_chanX_n3_driver_mux_fanins  <= "0" & CLB_8_1_OUT_pin_2 & track_8_1_chanY_n8 & track_8_2_chanY_n9;
	track_8_1_chanX_n4_driver_mux_fanins  <= CLB_8_1_OUT_pin_2 & track_7_1_chanY_n8 & track_7_1_chanX_n4 & track_7_2_chanY_n3;
	track_8_1_chanX_n5_driver_mux_fanins  <= "0" & CLB_8_1_OUT_pin_2 & track_8_1_chanY_n10 & track_8_2_chanY_n11;
	track_8_1_chanX_n6_driver_mux_fanins  <= CLB_8_1_OUT_pin_2 & track_7_1_chanY_n6 & track_7_1_chanX_n6 & track_7_2_chanY_n5;
	track_8_1_chanX_n7_driver_mux_fanins  <= "0" & CLB_8_1_OUT_pin_2 & track_8_1_chanY_n12 & track_8_2_chanY_n13;
	track_8_1_chanX_n8_driver_mux_fanins  <= CLB_8_2_OUT_pin_0 & track_7_1_chanY_n4 & track_7_1_chanX_n8 & track_7_2_chanY_n7;
	track_8_1_chanX_n9_driver_mux_fanins  <= "0" & CLB_8_2_OUT_pin_0 & track_8_1_chanY_n2 & track_8_2_chanY_n3;
	track_8_1_chanY_n0_driver_mux_fanins  <= "0" & IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_0_chanX_n0;
	track_8_1_chanY_n1_driver_mux_fanins  <= IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_1_chanX_n0 & track_8_2_chanY_n1;
	track_8_1_chanY_n10_driver_mux_fanins <= IO_9_1_OUT_pin_0 & track_8_0_chanX_n6;
	track_8_1_chanY_n11_driver_mux_fanins <= "0" & IO_9_1_OUT_pin_0 & track_8_1_chanX_n10 & track_8_2_chanY_n11;
	track_8_1_chanY_n12_driver_mux_fanins <= IO_9_1_OUT_pin_0 & track_8_0_chanX_n4;
	track_8_1_chanY_n13_driver_mux_fanins <= "0" & IO_9_1_OUT_pin_0 & track_8_1_chanX_n12 & track_8_2_chanY_n13;
	track_8_1_chanY_n14_driver_mux_fanins <= IO_9_1_OUT_pin_0 & track_8_0_chanX_n2;
	track_8_1_chanY_n15_driver_mux_fanins <= "0" & IO_9_1_OUT_pin_0 & track_8_1_chanX_n14 & track_8_2_chanY_n15;
	track_8_1_chanY_n2_driver_mux_fanins  <= "0" & IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_0_chanX_n14;
	track_8_1_chanY_n3_driver_mux_fanins  <= IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_1_chanX_n2 & track_8_2_chanY_n3;
	track_8_1_chanY_n4_driver_mux_fanins  <= "0" & IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_0_chanX_n12;
	track_8_1_chanY_n5_driver_mux_fanins  <= IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_1_chanX_n4 & track_8_2_chanY_n5;
	track_8_1_chanY_n6_driver_mux_fanins  <= "0" & IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_0_chanX_n10;
	track_8_1_chanY_n7_driver_mux_fanins  <= IO_9_1_OUT_pin_1 & CLB_8_1_OUT_pin_3 & track_8_1_chanX_n6 & track_8_2_chanY_n7;
	track_8_1_chanY_n8_driver_mux_fanins  <= IO_9_1_OUT_pin_0 & track_8_0_chanX_n8;
	track_8_1_chanY_n9_driver_mux_fanins  <= "0" & IO_9_1_OUT_pin_0 & track_8_1_chanX_n8 & track_8_2_chanY_n9;
	track_8_2_chanX_n0_driver_mux_fanins  <= CLB_8_2_OUT_pin_2 & track_7_2_chanY_n12 & track_7_2_chanX_n0 & track_7_3_chanY_n15;
	track_8_2_chanX_n1_driver_mux_fanins  <= "0" & CLB_8_2_OUT_pin_2 & track_8_2_chanY_n0 & track_8_3_chanY_n1;
	track_8_2_chanX_n10_driver_mux_fanins <= CLB_8_3_OUT_pin_0 & track_7_2_chanY_n2 & track_7_2_chanX_n10 & track_7_3_chanY_n9;
	track_8_2_chanX_n11_driver_mux_fanins <= "0" & CLB_8_3_OUT_pin_0 & track_8_2_chanY_n4 & track_8_3_chanY_n5;
	track_8_2_chanX_n12_driver_mux_fanins <= CLB_8_3_OUT_pin_0 & track_7_2_chanY_n0 & track_7_2_chanX_n12 & track_7_3_chanY_n11;
	track_8_2_chanX_n13_driver_mux_fanins <= "0" & CLB_8_3_OUT_pin_0 & track_8_2_chanY_n6 & track_8_3_chanY_n7;
	track_8_2_chanX_n14_driver_mux_fanins <= CLB_8_3_OUT_pin_0 & track_7_2_chanY_n14 & track_7_2_chanX_n14 & track_7_3_chanY_n13;
	track_8_2_chanX_n15_driver_mux_fanins <= "0" & CLB_8_3_OUT_pin_0 & track_8_2_chanY_n14 & track_8_3_chanY_n15;
	track_8_2_chanX_n2_driver_mux_fanins  <= CLB_8_2_OUT_pin_2 & track_7_2_chanY_n10 & track_7_2_chanX_n2 & track_7_3_chanY_n1;
	track_8_2_chanX_n3_driver_mux_fanins  <= "0" & CLB_8_2_OUT_pin_2 & track_8_2_chanY_n8 & track_8_3_chanY_n9;
	track_8_2_chanX_n4_driver_mux_fanins  <= CLB_8_2_OUT_pin_2 & track_7_2_chanY_n8 & track_7_2_chanX_n4 & track_7_3_chanY_n3;
	track_8_2_chanX_n5_driver_mux_fanins  <= "0" & CLB_8_2_OUT_pin_2 & track_8_2_chanY_n10 & track_8_3_chanY_n11;
	track_8_2_chanX_n6_driver_mux_fanins  <= CLB_8_2_OUT_pin_2 & track_7_2_chanY_n6 & track_7_2_chanX_n6 & track_7_3_chanY_n5;
	track_8_2_chanX_n7_driver_mux_fanins  <= "0" & CLB_8_2_OUT_pin_2 & track_8_2_chanY_n12 & track_8_3_chanY_n13;
	track_8_2_chanX_n8_driver_mux_fanins  <= CLB_8_3_OUT_pin_0 & track_7_2_chanY_n4 & track_7_2_chanX_n8 & track_7_3_chanY_n7;
	track_8_2_chanX_n9_driver_mux_fanins  <= "0" & CLB_8_3_OUT_pin_0 & track_8_2_chanY_n2 & track_8_3_chanY_n3;
	track_8_2_chanY_n0_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_1_chanY_n0 & track_8_1_chanX_n0;
	track_8_2_chanY_n1_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_2_chanX_n0 & track_8_3_chanY_n1;
	track_8_2_chanY_n10_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_1_chanY_n10 & track_8_1_chanX_n10;
	track_8_2_chanY_n11_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_2_chanX_n10 & track_8_3_chanY_n11;
	track_8_2_chanY_n12_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_1_chanY_n12 & track_8_1_chanX_n12;
	track_8_2_chanY_n13_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_2_chanX_n12 & track_8_3_chanY_n13;
	track_8_2_chanY_n14_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_1_chanY_n14 & track_8_1_chanX_n14;
	track_8_2_chanY_n15_driver_mux_fanins <= "0" & IO_9_2_OUT_pin_0 & track_8_2_chanX_n14 & track_8_3_chanY_n15;
	track_8_2_chanY_n2_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_1_chanY_n2 & track_8_1_chanX_n2;
	track_8_2_chanY_n3_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_2_chanX_n2 & track_8_3_chanY_n3;
	track_8_2_chanY_n4_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_1_chanY_n4 & track_8_1_chanX_n4;
	track_8_2_chanY_n5_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_2_chanX_n4 & track_8_3_chanY_n5;
	track_8_2_chanY_n6_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_1_chanY_n6 & track_8_1_chanX_n6;
	track_8_2_chanY_n7_driver_mux_fanins  <= IO_9_2_OUT_pin_1 & CLB_8_2_OUT_pin_3 & track_8_2_chanX_n6 & track_8_3_chanY_n7;
	track_8_2_chanY_n8_driver_mux_fanins  <= "0" & IO_9_2_OUT_pin_0 & track_8_1_chanY_n8 & track_8_1_chanX_n8;
	track_8_2_chanY_n9_driver_mux_fanins  <= "0" & IO_9_2_OUT_pin_0 & track_8_2_chanX_n8 & track_8_3_chanY_n9;
	track_8_3_chanX_n0_driver_mux_fanins  <= CLB_8_3_OUT_pin_2 & track_7_3_chanY_n12 & track_7_3_chanX_n0 & track_7_4_chanY_n15;
	track_8_3_chanX_n1_driver_mux_fanins  <= "0" & CLB_8_3_OUT_pin_2 & track_8_3_chanY_n0 & track_8_4_chanY_n1;
	track_8_3_chanX_n10_driver_mux_fanins <= CLB_8_4_OUT_pin_0 & track_7_3_chanY_n2 & track_7_3_chanX_n10 & track_7_4_chanY_n9;
	track_8_3_chanX_n11_driver_mux_fanins <= "0" & CLB_8_4_OUT_pin_0 & track_8_3_chanY_n4 & track_8_4_chanY_n5;
	track_8_3_chanX_n12_driver_mux_fanins <= CLB_8_4_OUT_pin_0 & track_7_3_chanY_n0 & track_7_3_chanX_n12 & track_7_4_chanY_n11;
	track_8_3_chanX_n13_driver_mux_fanins <= "0" & CLB_8_4_OUT_pin_0 & track_8_3_chanY_n6 & track_8_4_chanY_n7;
	track_8_3_chanX_n14_driver_mux_fanins <= CLB_8_4_OUT_pin_0 & track_7_3_chanY_n14 & track_7_3_chanX_n14 & track_7_4_chanY_n13;
	track_8_3_chanX_n15_driver_mux_fanins <= "0" & CLB_8_4_OUT_pin_0 & track_8_3_chanY_n14 & track_8_4_chanY_n15;
	track_8_3_chanX_n2_driver_mux_fanins  <= CLB_8_3_OUT_pin_2 & track_7_3_chanY_n10 & track_7_3_chanX_n2 & track_7_4_chanY_n1;
	track_8_3_chanX_n3_driver_mux_fanins  <= "0" & CLB_8_3_OUT_pin_2 & track_8_3_chanY_n8 & track_8_4_chanY_n9;
	track_8_3_chanX_n4_driver_mux_fanins  <= CLB_8_3_OUT_pin_2 & track_7_3_chanY_n8 & track_7_3_chanX_n4 & track_7_4_chanY_n3;
	track_8_3_chanX_n5_driver_mux_fanins  <= "0" & CLB_8_3_OUT_pin_2 & track_8_3_chanY_n10 & track_8_4_chanY_n11;
	track_8_3_chanX_n6_driver_mux_fanins  <= CLB_8_3_OUT_pin_2 & track_7_3_chanY_n6 & track_7_3_chanX_n6 & track_7_4_chanY_n5;
	track_8_3_chanX_n7_driver_mux_fanins  <= "0" & CLB_8_3_OUT_pin_2 & track_8_3_chanY_n12 & track_8_4_chanY_n13;
	track_8_3_chanX_n8_driver_mux_fanins  <= CLB_8_4_OUT_pin_0 & track_7_3_chanY_n4 & track_7_3_chanX_n8 & track_7_4_chanY_n7;
	track_8_3_chanX_n9_driver_mux_fanins  <= "0" & CLB_8_4_OUT_pin_0 & track_8_3_chanY_n2 & track_8_4_chanY_n3;
	track_8_3_chanY_n0_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_2_chanY_n0 & track_8_2_chanX_n0;
	track_8_3_chanY_n1_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_3_chanX_n0 & track_8_4_chanY_n1;
	track_8_3_chanY_n10_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_2_chanY_n10 & track_8_2_chanX_n10;
	track_8_3_chanY_n11_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_3_chanX_n10 & track_8_4_chanY_n11;
	track_8_3_chanY_n12_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_2_chanY_n12 & track_8_2_chanX_n12;
	track_8_3_chanY_n13_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_3_chanX_n12 & track_8_4_chanY_n13;
	track_8_3_chanY_n14_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_2_chanY_n14 & track_8_2_chanX_n14;
	track_8_3_chanY_n15_driver_mux_fanins <= "0" & IO_9_3_OUT_pin_0 & track_8_3_chanX_n14 & track_8_4_chanY_n15;
	track_8_3_chanY_n2_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_2_chanY_n2 & track_8_2_chanX_n2;
	track_8_3_chanY_n3_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_3_chanX_n2 & track_8_4_chanY_n3;
	track_8_3_chanY_n4_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_2_chanY_n4 & track_8_2_chanX_n4;
	track_8_3_chanY_n5_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_3_chanX_n4 & track_8_4_chanY_n5;
	track_8_3_chanY_n6_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_2_chanY_n6 & track_8_2_chanX_n6;
	track_8_3_chanY_n7_driver_mux_fanins  <= IO_9_3_OUT_pin_1 & CLB_8_3_OUT_pin_3 & track_8_3_chanX_n6 & track_8_4_chanY_n7;
	track_8_3_chanY_n8_driver_mux_fanins  <= "0" & IO_9_3_OUT_pin_0 & track_8_2_chanY_n8 & track_8_2_chanX_n8;
	track_8_3_chanY_n9_driver_mux_fanins  <= "0" & IO_9_3_OUT_pin_0 & track_8_3_chanX_n8 & track_8_4_chanY_n9;
	track_8_4_chanX_n0_driver_mux_fanins  <= CLB_8_4_OUT_pin_2 & track_7_4_chanY_n12 & track_7_4_chanX_n0 & track_7_5_chanY_n15;
	track_8_4_chanX_n1_driver_mux_fanins  <= "0" & CLB_8_4_OUT_pin_2 & track_8_4_chanY_n0 & track_8_5_chanY_n1;
	track_8_4_chanX_n10_driver_mux_fanins <= CLB_8_5_OUT_pin_0 & track_7_4_chanY_n2 & track_7_4_chanX_n10 & track_7_5_chanY_n9;
	track_8_4_chanX_n11_driver_mux_fanins <= "0" & CLB_8_5_OUT_pin_0 & track_8_4_chanY_n4 & track_8_5_chanY_n5;
	track_8_4_chanX_n12_driver_mux_fanins <= CLB_8_5_OUT_pin_0 & track_7_4_chanY_n0 & track_7_4_chanX_n12 & track_7_5_chanY_n11;
	track_8_4_chanX_n13_driver_mux_fanins <= "0" & CLB_8_5_OUT_pin_0 & track_8_4_chanY_n6 & track_8_5_chanY_n7;
	track_8_4_chanX_n14_driver_mux_fanins <= CLB_8_5_OUT_pin_0 & track_7_4_chanY_n14 & track_7_4_chanX_n14 & track_7_5_chanY_n13;
	track_8_4_chanX_n15_driver_mux_fanins <= "0" & CLB_8_5_OUT_pin_0 & track_8_4_chanY_n14 & track_8_5_chanY_n15;
	track_8_4_chanX_n2_driver_mux_fanins  <= CLB_8_4_OUT_pin_2 & track_7_4_chanY_n10 & track_7_4_chanX_n2 & track_7_5_chanY_n1;
	track_8_4_chanX_n3_driver_mux_fanins  <= "0" & CLB_8_4_OUT_pin_2 & track_8_4_chanY_n8 & track_8_5_chanY_n9;
	track_8_4_chanX_n4_driver_mux_fanins  <= CLB_8_4_OUT_pin_2 & track_7_4_chanY_n8 & track_7_4_chanX_n4 & track_7_5_chanY_n3;
	track_8_4_chanX_n5_driver_mux_fanins  <= "0" & CLB_8_4_OUT_pin_2 & track_8_4_chanY_n10 & track_8_5_chanY_n11;
	track_8_4_chanX_n6_driver_mux_fanins  <= CLB_8_4_OUT_pin_2 & track_7_4_chanY_n6 & track_7_4_chanX_n6 & track_7_5_chanY_n5;
	track_8_4_chanX_n7_driver_mux_fanins  <= "0" & CLB_8_4_OUT_pin_2 & track_8_4_chanY_n12 & track_8_5_chanY_n13;
	track_8_4_chanX_n8_driver_mux_fanins  <= CLB_8_5_OUT_pin_0 & track_7_4_chanY_n4 & track_7_4_chanX_n8 & track_7_5_chanY_n7;
	track_8_4_chanX_n9_driver_mux_fanins  <= "0" & CLB_8_5_OUT_pin_0 & track_8_4_chanY_n2 & track_8_5_chanY_n3;
	track_8_4_chanY_n0_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_3_chanY_n0 & track_8_3_chanX_n0;
	track_8_4_chanY_n1_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_4_chanX_n0 & track_8_5_chanY_n1;
	track_8_4_chanY_n10_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_3_chanY_n10 & track_8_3_chanX_n10;
	track_8_4_chanY_n11_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_4_chanX_n10 & track_8_5_chanY_n11;
	track_8_4_chanY_n12_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_3_chanY_n12 & track_8_3_chanX_n12;
	track_8_4_chanY_n13_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_4_chanX_n12 & track_8_5_chanY_n13;
	track_8_4_chanY_n14_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_3_chanY_n14 & track_8_3_chanX_n14;
	track_8_4_chanY_n15_driver_mux_fanins <= "0" & IO_9_4_OUT_pin_0 & track_8_4_chanX_n14 & track_8_5_chanY_n15;
	track_8_4_chanY_n2_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_3_chanY_n2 & track_8_3_chanX_n2;
	track_8_4_chanY_n3_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_4_chanX_n2 & track_8_5_chanY_n3;
	track_8_4_chanY_n4_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_3_chanY_n4 & track_8_3_chanX_n4;
	track_8_4_chanY_n5_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_4_chanX_n4 & track_8_5_chanY_n5;
	track_8_4_chanY_n6_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_3_chanY_n6 & track_8_3_chanX_n6;
	track_8_4_chanY_n7_driver_mux_fanins  <= IO_9_4_OUT_pin_1 & CLB_8_4_OUT_pin_3 & track_8_4_chanX_n6 & track_8_5_chanY_n7;
	track_8_4_chanY_n8_driver_mux_fanins  <= "0" & IO_9_4_OUT_pin_0 & track_8_3_chanY_n8 & track_8_3_chanX_n8;
	track_8_4_chanY_n9_driver_mux_fanins  <= "0" & IO_9_4_OUT_pin_0 & track_8_4_chanX_n8 & track_8_5_chanY_n9;
	track_8_5_chanX_n0_driver_mux_fanins  <= CLB_8_5_OUT_pin_2 & track_7_5_chanY_n12 & track_7_5_chanX_n0 & track_7_6_chanY_n15;
	track_8_5_chanX_n1_driver_mux_fanins  <= "0" & CLB_8_5_OUT_pin_2 & track_8_5_chanY_n0 & track_8_6_chanY_n1;
	track_8_5_chanX_n10_driver_mux_fanins <= CLB_8_6_OUT_pin_0 & track_7_5_chanY_n2 & track_7_5_chanX_n10 & track_7_6_chanY_n9;
	track_8_5_chanX_n11_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_0 & track_8_5_chanY_n4 & track_8_6_chanY_n5;
	track_8_5_chanX_n12_driver_mux_fanins <= CLB_8_6_OUT_pin_0 & track_7_5_chanY_n0 & track_7_5_chanX_n12 & track_7_6_chanY_n11;
	track_8_5_chanX_n13_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_0 & track_8_5_chanY_n6 & track_8_6_chanY_n7;
	track_8_5_chanX_n14_driver_mux_fanins <= CLB_8_6_OUT_pin_0 & track_7_5_chanY_n14 & track_7_5_chanX_n14 & track_7_6_chanY_n13;
	track_8_5_chanX_n15_driver_mux_fanins <= "0" & CLB_8_6_OUT_pin_0 & track_8_5_chanY_n14 & track_8_6_chanY_n15;
	track_8_5_chanX_n2_driver_mux_fanins  <= CLB_8_5_OUT_pin_2 & track_7_5_chanY_n10 & track_7_5_chanX_n2 & track_7_6_chanY_n1;
	track_8_5_chanX_n3_driver_mux_fanins  <= "0" & CLB_8_5_OUT_pin_2 & track_8_5_chanY_n8 & track_8_6_chanY_n9;
	track_8_5_chanX_n4_driver_mux_fanins  <= CLB_8_5_OUT_pin_2 & track_7_5_chanY_n8 & track_7_5_chanX_n4 & track_7_6_chanY_n3;
	track_8_5_chanX_n5_driver_mux_fanins  <= "0" & CLB_8_5_OUT_pin_2 & track_8_5_chanY_n10 & track_8_6_chanY_n11;
	track_8_5_chanX_n6_driver_mux_fanins  <= CLB_8_5_OUT_pin_2 & track_7_5_chanY_n6 & track_7_5_chanX_n6 & track_7_6_chanY_n5;
	track_8_5_chanX_n7_driver_mux_fanins  <= "0" & CLB_8_5_OUT_pin_2 & track_8_5_chanY_n12 & track_8_6_chanY_n13;
	track_8_5_chanX_n8_driver_mux_fanins  <= CLB_8_6_OUT_pin_0 & track_7_5_chanY_n4 & track_7_5_chanX_n8 & track_7_6_chanY_n7;
	track_8_5_chanX_n9_driver_mux_fanins  <= "0" & CLB_8_6_OUT_pin_0 & track_8_5_chanY_n2 & track_8_6_chanY_n3;
	track_8_5_chanY_n0_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_4_chanY_n0 & track_8_4_chanX_n0;
	track_8_5_chanY_n1_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_5_chanX_n0 & track_8_6_chanY_n1;
	track_8_5_chanY_n10_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_4_chanY_n10 & track_8_4_chanX_n10;
	track_8_5_chanY_n11_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_5_chanX_n10 & track_8_6_chanY_n11;
	track_8_5_chanY_n12_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_4_chanY_n12 & track_8_4_chanX_n12;
	track_8_5_chanY_n13_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_5_chanX_n12 & track_8_6_chanY_n13;
	track_8_5_chanY_n14_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_4_chanY_n14 & track_8_4_chanX_n14;
	track_8_5_chanY_n15_driver_mux_fanins <= "0" & IO_9_5_OUT_pin_0 & track_8_5_chanX_n14 & track_8_6_chanY_n15;
	track_8_5_chanY_n2_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_4_chanY_n2 & track_8_4_chanX_n2;
	track_8_5_chanY_n3_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_5_chanX_n2 & track_8_6_chanY_n3;
	track_8_5_chanY_n4_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_4_chanY_n4 & track_8_4_chanX_n4;
	track_8_5_chanY_n5_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_5_chanX_n4 & track_8_6_chanY_n5;
	track_8_5_chanY_n6_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_4_chanY_n6 & track_8_4_chanX_n6;
	track_8_5_chanY_n7_driver_mux_fanins  <= IO_9_5_OUT_pin_1 & CLB_8_5_OUT_pin_3 & track_8_5_chanX_n6 & track_8_6_chanY_n7;
	track_8_5_chanY_n8_driver_mux_fanins  <= "0" & IO_9_5_OUT_pin_0 & track_8_4_chanY_n8 & track_8_4_chanX_n8;
	track_8_5_chanY_n9_driver_mux_fanins  <= "0" & IO_9_5_OUT_pin_0 & track_8_5_chanX_n8 & track_8_6_chanY_n9;
	track_8_6_chanX_n0_driver_mux_fanins  <= IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_7_6_chanY_n0 & track_7_6_chanX_n0;
	track_8_6_chanX_n1_driver_mux_fanins  <= "0" & IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_8_6_chanY_n14;
	track_8_6_chanX_n10_driver_mux_fanins <= "0" & IO_8_7_OUT_pin_0 & track_7_6_chanY_n10 & track_7_6_chanX_n10;
	track_8_6_chanX_n11_driver_mux_fanins <= IO_8_7_OUT_pin_0 & track_8_6_chanY_n8;
	track_8_6_chanX_n12_driver_mux_fanins <= "0" & IO_8_7_OUT_pin_0 & track_7_6_chanY_n12 & track_7_6_chanX_n12;
	track_8_6_chanX_n13_driver_mux_fanins <= IO_8_7_OUT_pin_0 & track_8_6_chanY_n10;
	track_8_6_chanX_n14_driver_mux_fanins <= "0" & IO_8_7_OUT_pin_0 & track_7_6_chanY_n14 & track_7_6_chanX_n14;
	track_8_6_chanX_n15_driver_mux_fanins <= IO_8_7_OUT_pin_0 & track_8_6_chanY_n12;
	track_8_6_chanX_n2_driver_mux_fanins  <= IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_7_6_chanY_n2 & track_7_6_chanX_n2;
	track_8_6_chanX_n3_driver_mux_fanins  <= "0" & IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_8_6_chanY_n0;
	track_8_6_chanX_n4_driver_mux_fanins  <= IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_7_6_chanY_n4 & track_7_6_chanX_n4;
	track_8_6_chanX_n5_driver_mux_fanins  <= "0" & IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_8_6_chanY_n2;
	track_8_6_chanX_n6_driver_mux_fanins  <= IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_7_6_chanY_n6 & track_7_6_chanX_n6;
	track_8_6_chanX_n7_driver_mux_fanins  <= "0" & IO_8_7_OUT_pin_1 & CLB_8_6_OUT_pin_2 & track_8_6_chanY_n4;
	track_8_6_chanX_n8_driver_mux_fanins  <= "0" & IO_8_7_OUT_pin_0 & track_7_6_chanY_n8 & track_7_6_chanX_n8;
	track_8_6_chanX_n9_driver_mux_fanins  <= IO_8_7_OUT_pin_0 & track_8_6_chanY_n6;
	track_8_6_chanY_n0_driver_mux_fanins  <= IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_5_chanY_n0 & track_8_5_chanX_n0;
	track_8_6_chanY_n1_driver_mux_fanins  <= "0" & IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_6_chanX_n2;
	track_8_6_chanY_n10_driver_mux_fanins <= "0" & IO_9_6_OUT_pin_0 & track_8_5_chanY_n10 & track_8_5_chanX_n10;
	track_8_6_chanY_n11_driver_mux_fanins <= IO_9_6_OUT_pin_0 & track_8_6_chanX_n12;
	track_8_6_chanY_n12_driver_mux_fanins <= "0" & IO_9_6_OUT_pin_0 & track_8_5_chanY_n12 & track_8_5_chanX_n12;
	track_8_6_chanY_n13_driver_mux_fanins <= IO_9_6_OUT_pin_0 & track_8_6_chanX_n14;
	track_8_6_chanY_n14_driver_mux_fanins <= "0" & IO_9_6_OUT_pin_0 & track_8_5_chanY_n14 & track_8_5_chanX_n14;
	track_8_6_chanY_n15_driver_mux_fanins <= IO_9_6_OUT_pin_0 & track_8_6_chanX_n0;
	track_8_6_chanY_n2_driver_mux_fanins  <= IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_5_chanY_n2 & track_8_5_chanX_n2;
	track_8_6_chanY_n3_driver_mux_fanins  <= "0" & IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_6_chanX_n4;
	track_8_6_chanY_n4_driver_mux_fanins  <= IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_5_chanY_n4 & track_8_5_chanX_n4;
	track_8_6_chanY_n5_driver_mux_fanins  <= "0" & IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_6_chanX_n6;
	track_8_6_chanY_n6_driver_mux_fanins  <= IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_5_chanY_n6 & track_8_5_chanX_n6;
	track_8_6_chanY_n7_driver_mux_fanins  <= "0" & IO_9_6_OUT_pin_1 & CLB_8_6_OUT_pin_3 & track_8_6_chanX_n8;
	track_8_6_chanY_n8_driver_mux_fanins  <= "0" & IO_9_6_OUT_pin_0 & track_8_5_chanY_n8 & track_8_5_chanX_n8;
	track_8_6_chanY_n9_driver_mux_fanins  <= IO_9_6_OUT_pin_0 & track_8_6_chanX_n10;

	-- Tracks selectors (selector of the mux driving the track, i.e. the bitstream portion configuring the track) --
	track_0_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7465 downto 7464)));
	track_0_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7467 downto 7466)));
	track_0_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7468 downto 7468)));
	track_0_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7470 downto 7469)));
	track_0_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7471 downto 7471)));
	track_0_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7473 downto 7472)));
	track_0_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7474 downto 7474)));
	track_0_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7476 downto 7475)));
	track_0_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7478 downto 7477)));
	track_0_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7480 downto 7479)));
	track_0_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7482 downto 7481)));
	track_0_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7484 downto 7483)));
	track_0_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7486 downto 7485)));
	track_0_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7488 downto 7487)));
	track_0_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7489 downto 7489)));
	track_0_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7491 downto 7490)));
	track_0_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7493 downto 7492)));
	track_0_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7495 downto 7494)));
	track_0_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7497 downto 7496)));
	track_0_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7499 downto 7498)));
	track_0_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7501 downto 7500)));
	track_0_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7503 downto 7502)));
	track_0_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7505 downto 7504)));
	track_0_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7507 downto 7506)));
	track_0_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7509 downto 7508)));
	track_0_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7511 downto 7510)));
	track_0_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7513 downto 7512)));
	track_0_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7515 downto 7514)));
	track_0_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7517 downto 7516)));
	track_0_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7519 downto 7518)));
	track_0_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7521 downto 7520)));
	track_0_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7523 downto 7522)));
	track_0_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7525 downto 7524)));
	track_0_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7527 downto 7526)));
	track_0_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7529 downto 7528)));
	track_0_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7531 downto 7530)));
	track_0_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7533 downto 7532)));
	track_0_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7535 downto 7534)));
	track_0_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7537 downto 7536)));
	track_0_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7539 downto 7538)));
	track_0_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7541 downto 7540)));
	track_0_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7543 downto 7542)));
	track_0_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7545 downto 7544)));
	track_0_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7547 downto 7546)));
	track_0_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7549 downto 7548)));
	track_0_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7551 downto 7550)));
	track_0_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7553 downto 7552)));
	track_0_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7555 downto 7554)));
	track_0_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7557 downto 7556)));
	track_0_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7559 downto 7558)));
	track_0_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7561 downto 7560)));
	track_0_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7563 downto 7562)));
	track_0_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7565 downto 7564)));
	track_0_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7567 downto 7566)));
	track_0_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7569 downto 7568)));
	track_0_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7571 downto 7570)));
	track_0_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7573 downto 7572)));
	track_0_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7575 downto 7574)));
	track_0_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7577 downto 7576)));
	track_0_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7579 downto 7578)));
	track_0_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7581 downto 7580)));
	track_0_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7583 downto 7582)));
	track_0_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7585 downto 7584)));
	track_0_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7587 downto 7586)));
	track_0_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7589 downto 7588)));
	track_0_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7591 downto 7590)));
	track_0_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7593 downto 7592)));
	track_0_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7595 downto 7594)));
	track_0_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7597 downto 7596)));
	track_0_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7599 downto 7598)));
	track_0_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7601 downto 7600)));
	track_0_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7603 downto 7602)));
	track_0_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7605 downto 7604)));
	track_0_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7607 downto 7606)));
	track_0_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7609 downto 7608)));
	track_0_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7611 downto 7610)));
	track_0_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7613 downto 7612)));
	track_0_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7615 downto 7614)));
	track_0_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7617 downto 7616)));
	track_0_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7619 downto 7618)));
	track_0_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7621 downto 7620)));
	track_0_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7623 downto 7622)));
	track_0_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7625 downto 7624)));
	track_0_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7626 downto 7626)));
	track_0_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7628 downto 7627)));
	track_0_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7629 downto 7629)));
	track_0_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7631 downto 7630)));
	track_0_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7632 downto 7632)));
	track_0_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7634 downto 7633)));
	track_0_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7636 downto 7635)));
	track_0_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7638 downto 7637)));
	track_0_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7640 downto 7639)));
	track_0_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7642 downto 7641)));
	track_0_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7644 downto 7643)));
	track_0_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7646 downto 7645)));
	track_0_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7647 downto 7647)));
	track_1_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7649 downto 7648)));
	track_1_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7651 downto 7650)));
	track_1_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7652 downto 7652)));
	track_1_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7654 downto 7653)));
	track_1_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7655 downto 7655)));
	track_1_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7657 downto 7656)));
	track_1_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7658 downto 7658)));
	track_1_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7660 downto 7659)));
	track_1_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7662 downto 7661)));
	track_1_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7664 downto 7663)));
	track_1_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7666 downto 7665)));
	track_1_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7668 downto 7667)));
	track_1_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7670 downto 7669)));
	track_1_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7672 downto 7671)));
	track_1_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7673 downto 7673)));
	track_1_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7675 downto 7674)));
	track_1_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7677 downto 7676)));
	track_1_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7679 downto 7678)));
	track_1_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7681 downto 7680)));
	track_1_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7683 downto 7682)));
	track_1_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7685 downto 7684)));
	track_1_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7687 downto 7686)));
	track_1_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7689 downto 7688)));
	track_1_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7691 downto 7690)));
	track_1_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7693 downto 7692)));
	track_1_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7695 downto 7694)));
	track_1_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7697 downto 7696)));
	track_1_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7699 downto 7698)));
	track_1_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7701 downto 7700)));
	track_1_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7703 downto 7702)));
	track_1_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7705 downto 7704)));
	track_1_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7707 downto 7706)));
	track_1_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7709 downto 7708)));
	track_1_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7711 downto 7710)));
	track_1_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7713 downto 7712)));
	track_1_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7715 downto 7714)));
	track_1_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7717 downto 7716)));
	track_1_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7719 downto 7718)));
	track_1_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7721 downto 7720)));
	track_1_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7723 downto 7722)));
	track_1_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7725 downto 7724)));
	track_1_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7727 downto 7726)));
	track_1_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7729 downto 7728)));
	track_1_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7731 downto 7730)));
	track_1_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7733 downto 7732)));
	track_1_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7735 downto 7734)));
	track_1_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7737 downto 7736)));
	track_1_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7739 downto 7738)));
	track_1_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7741 downto 7740)));
	track_1_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7743 downto 7742)));
	track_1_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7745 downto 7744)));
	track_1_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7747 downto 7746)));
	track_1_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7749 downto 7748)));
	track_1_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7751 downto 7750)));
	track_1_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7753 downto 7752)));
	track_1_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7755 downto 7754)));
	track_1_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7757 downto 7756)));
	track_1_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7759 downto 7758)));
	track_1_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7761 downto 7760)));
	track_1_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7763 downto 7762)));
	track_1_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7765 downto 7764)));
	track_1_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7767 downto 7766)));
	track_1_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7769 downto 7768)));
	track_1_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7771 downto 7770)));
	track_1_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7773 downto 7772)));
	track_1_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7775 downto 7774)));
	track_1_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7777 downto 7776)));
	track_1_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7779 downto 7778)));
	track_1_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7781 downto 7780)));
	track_1_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7783 downto 7782)));
	track_1_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7785 downto 7784)));
	track_1_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7787 downto 7786)));
	track_1_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7789 downto 7788)));
	track_1_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7791 downto 7790)));
	track_1_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7793 downto 7792)));
	track_1_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7795 downto 7794)));
	track_1_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7797 downto 7796)));
	track_1_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7799 downto 7798)));
	track_1_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7801 downto 7800)));
	track_1_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7803 downto 7802)));
	track_1_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7805 downto 7804)));
	track_1_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7807 downto 7806)));
	track_1_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7809 downto 7808)));
	track_1_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7811 downto 7810)));
	track_1_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7813 downto 7812)));
	track_1_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7815 downto 7814)));
	track_1_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7817 downto 7816)));
	track_1_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7819 downto 7818)));
	track_1_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7821 downto 7820)));
	track_1_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7823 downto 7822)));
	track_1_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7825 downto 7824)));
	track_1_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7827 downto 7826)));
	track_1_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7829 downto 7828)));
	track_1_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7831 downto 7830)));
	track_1_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7833 downto 7832)));
	track_1_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7835 downto 7834)));
	track_1_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7837 downto 7836)));
	track_1_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7839 downto 7838)));
	track_1_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7841 downto 7840)));
	track_1_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7843 downto 7842)));
	track_1_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7845 downto 7844)));
	track_1_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7847 downto 7846)));
	track_1_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7849 downto 7848)));
	track_1_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7851 downto 7850)));
	track_1_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7853 downto 7852)));
	track_1_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7855 downto 7854)));
	track_1_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7857 downto 7856)));
	track_1_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7859 downto 7858)));
	track_1_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7861 downto 7860)));
	track_1_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7863 downto 7862)));
	track_1_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7865 downto 7864)));
	track_1_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7867 downto 7866)));
	track_1_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7869 downto 7868)));
	track_1_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7871 downto 7870)));
	track_1_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7873 downto 7872)));
	track_1_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7875 downto 7874)));
	track_1_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7877 downto 7876)));
	track_1_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7879 downto 7878)));
	track_1_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7881 downto 7880)));
	track_1_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7883 downto 7882)));
	track_1_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7885 downto 7884)));
	track_1_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7887 downto 7886)));
	track_1_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7889 downto 7888)));
	track_1_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7891 downto 7890)));
	track_1_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7893 downto 7892)));
	track_1_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7895 downto 7894)));
	track_1_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7897 downto 7896)));
	track_1_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7899 downto 7898)));
	track_1_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7901 downto 7900)));
	track_1_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7903 downto 7902)));
	track_1_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7905 downto 7904)));
	track_1_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7907 downto 7906)));
	track_1_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7909 downto 7908)));
	track_1_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7911 downto 7910)));
	track_1_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7913 downto 7912)));
	track_1_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7915 downto 7914)));
	track_1_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7917 downto 7916)));
	track_1_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7919 downto 7918)));
	track_1_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7921 downto 7920)));
	track_1_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7923 downto 7922)));
	track_1_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7925 downto 7924)));
	track_1_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7927 downto 7926)));
	track_1_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7929 downto 7928)));
	track_1_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7931 downto 7930)));
	track_1_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7933 downto 7932)));
	track_1_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7935 downto 7934)));
	track_1_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(7937 downto 7936)));
	track_1_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(7939 downto 7938)));
	track_1_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(7941 downto 7940)));
	track_1_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(7943 downto 7942)));
	track_1_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(7945 downto 7944)));
	track_1_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(7947 downto 7946)));
	track_1_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(7949 downto 7948)));
	track_1_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(7951 downto 7950)));
	track_1_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(7953 downto 7952)));
	track_1_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(7955 downto 7954)));
	track_1_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(7957 downto 7956)));
	track_1_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(7959 downto 7958)));
	track_1_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(7961 downto 7960)));
	track_1_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(7963 downto 7962)));
	track_1_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(7965 downto 7964)));
	track_1_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(7967 downto 7966)));
	track_1_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(7969 downto 7968)));
	track_1_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(7971 downto 7970)));
	track_1_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(7973 downto 7972)));
	track_1_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(7975 downto 7974)));
	track_1_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(7977 downto 7976)));
	track_1_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(7979 downto 7978)));
	track_1_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(7981 downto 7980)));
	track_1_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(7983 downto 7982)));
	track_1_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(7985 downto 7984)));
	track_1_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(7987 downto 7986)));
	track_1_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(7989 downto 7988)));
	track_1_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(7991 downto 7990)));
	track_1_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(7993 downto 7992)));
	track_1_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(7995 downto 7994)));
	track_1_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(7997 downto 7996)));
	track_1_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(7999 downto 7998)));
	track_1_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8000 downto 8000)));
	track_1_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8002 downto 8001)));
	track_1_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8003 downto 8003)));
	track_1_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8005 downto 8004)));
	track_1_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8006 downto 8006)));
	track_1_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8008 downto 8007)));
	track_1_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8010 downto 8009)));
	track_1_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8012 downto 8011)));
	track_1_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8014 downto 8013)));
	track_1_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8016 downto 8015)));
	track_1_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8018 downto 8017)));
	track_1_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8020 downto 8019)));
	track_1_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8021 downto 8021)));
	track_1_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8023 downto 8022)));
	track_1_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8025 downto 8024)));
	track_1_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8027 downto 8026)));
	track_1_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8029 downto 8028)));
	track_1_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8031 downto 8030)));
	track_1_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8033 downto 8032)));
	track_1_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8035 downto 8034)));
	track_1_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8037 downto 8036)));
	track_1_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8039 downto 8038)));
	track_1_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8041 downto 8040)));
	track_1_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8043 downto 8042)));
	track_1_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8045 downto 8044)));
	track_1_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8047 downto 8046)));
	track_1_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8049 downto 8048)));
	track_1_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8051 downto 8050)));
	track_1_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8053 downto 8052)));
	track_1_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8055 downto 8054)));
	track_2_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8057 downto 8056)));
	track_2_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8059 downto 8058)));
	track_2_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8061 downto 8060)));
	track_2_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8063 downto 8062)));
	track_2_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8065 downto 8064)));
	track_2_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8067 downto 8066)));
	track_2_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8069 downto 8068)));
	track_2_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8071 downto 8070)));
	track_2_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8073 downto 8072)));
	track_2_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8075 downto 8074)));
	track_2_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8077 downto 8076)));
	track_2_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8079 downto 8078)));
	track_2_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8081 downto 8080)));
	track_2_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8083 downto 8082)));
	track_2_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8085 downto 8084)));
	track_2_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8087 downto 8086)));
	track_2_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8089 downto 8088)));
	track_2_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8091 downto 8090)));
	track_2_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8093 downto 8092)));
	track_2_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8095 downto 8094)));
	track_2_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8097 downto 8096)));
	track_2_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8099 downto 8098)));
	track_2_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8101 downto 8100)));
	track_2_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8103 downto 8102)));
	track_2_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8105 downto 8104)));
	track_2_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8107 downto 8106)));
	track_2_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8109 downto 8108)));
	track_2_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8111 downto 8110)));
	track_2_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8113 downto 8112)));
	track_2_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8115 downto 8114)));
	track_2_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8117 downto 8116)));
	track_2_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8119 downto 8118)));
	track_2_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8121 downto 8120)));
	track_2_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8123 downto 8122)));
	track_2_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8125 downto 8124)));
	track_2_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8127 downto 8126)));
	track_2_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8129 downto 8128)));
	track_2_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8131 downto 8130)));
	track_2_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8133 downto 8132)));
	track_2_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8135 downto 8134)));
	track_2_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8137 downto 8136)));
	track_2_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8139 downto 8138)));
	track_2_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8141 downto 8140)));
	track_2_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8143 downto 8142)));
	track_2_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8145 downto 8144)));
	track_2_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8147 downto 8146)));
	track_2_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8149 downto 8148)));
	track_2_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8151 downto 8150)));
	track_2_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8153 downto 8152)));
	track_2_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8155 downto 8154)));
	track_2_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8157 downto 8156)));
	track_2_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8159 downto 8158)));
	track_2_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8161 downto 8160)));
	track_2_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8163 downto 8162)));
	track_2_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8165 downto 8164)));
	track_2_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8167 downto 8166)));
	track_2_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8169 downto 8168)));
	track_2_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8171 downto 8170)));
	track_2_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8173 downto 8172)));
	track_2_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8175 downto 8174)));
	track_2_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8177 downto 8176)));
	track_2_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8179 downto 8178)));
	track_2_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8181 downto 8180)));
	track_2_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8183 downto 8182)));
	track_2_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8185 downto 8184)));
	track_2_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8187 downto 8186)));
	track_2_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8189 downto 8188)));
	track_2_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8191 downto 8190)));
	track_2_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8193 downto 8192)));
	track_2_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8195 downto 8194)));
	track_2_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8197 downto 8196)));
	track_2_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8199 downto 8198)));
	track_2_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8201 downto 8200)));
	track_2_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8203 downto 8202)));
	track_2_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8205 downto 8204)));
	track_2_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8207 downto 8206)));
	track_2_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8209 downto 8208)));
	track_2_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8211 downto 8210)));
	track_2_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8213 downto 8212)));
	track_2_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8215 downto 8214)));
	track_2_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8217 downto 8216)));
	track_2_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8219 downto 8218)));
	track_2_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8221 downto 8220)));
	track_2_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8223 downto 8222)));
	track_2_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8225 downto 8224)));
	track_2_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8227 downto 8226)));
	track_2_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8229 downto 8228)));
	track_2_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8231 downto 8230)));
	track_2_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8233 downto 8232)));
	track_2_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8235 downto 8234)));
	track_2_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8237 downto 8236)));
	track_2_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8239 downto 8238)));
	track_2_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8241 downto 8240)));
	track_2_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8243 downto 8242)));
	track_2_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8245 downto 8244)));
	track_2_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8247 downto 8246)));
	track_2_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8249 downto 8248)));
	track_2_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8251 downto 8250)));
	track_2_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8253 downto 8252)));
	track_2_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8255 downto 8254)));
	track_2_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8257 downto 8256)));
	track_2_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8259 downto 8258)));
	track_2_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8261 downto 8260)));
	track_2_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8263 downto 8262)));
	track_2_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8265 downto 8264)));
	track_2_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8267 downto 8266)));
	track_2_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8269 downto 8268)));
	track_2_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8271 downto 8270)));
	track_2_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8273 downto 8272)));
	track_2_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8275 downto 8274)));
	track_2_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8277 downto 8276)));
	track_2_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8279 downto 8278)));
	track_2_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8281 downto 8280)));
	track_2_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8283 downto 8282)));
	track_2_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8285 downto 8284)));
	track_2_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8287 downto 8286)));
	track_2_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8289 downto 8288)));
	track_2_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8291 downto 8290)));
	track_2_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8293 downto 8292)));
	track_2_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8295 downto 8294)));
	track_2_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8297 downto 8296)));
	track_2_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8299 downto 8298)));
	track_2_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8301 downto 8300)));
	track_2_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8303 downto 8302)));
	track_2_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8305 downto 8304)));
	track_2_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8307 downto 8306)));
	track_2_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8309 downto 8308)));
	track_2_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8311 downto 8310)));
	track_2_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8313 downto 8312)));
	track_2_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8315 downto 8314)));
	track_2_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8317 downto 8316)));
	track_2_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8319 downto 8318)));
	track_2_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8321 downto 8320)));
	track_2_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8323 downto 8322)));
	track_2_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8325 downto 8324)));
	track_2_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8327 downto 8326)));
	track_2_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8329 downto 8328)));
	track_2_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8331 downto 8330)));
	track_2_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8333 downto 8332)));
	track_2_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8335 downto 8334)));
	track_2_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8337 downto 8336)));
	track_2_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8339 downto 8338)));
	track_2_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8341 downto 8340)));
	track_2_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8343 downto 8342)));
	track_2_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8345 downto 8344)));
	track_2_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8347 downto 8346)));
	track_2_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8349 downto 8348)));
	track_2_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8351 downto 8350)));
	track_2_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8353 downto 8352)));
	track_2_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8355 downto 8354)));
	track_2_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8357 downto 8356)));
	track_2_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8359 downto 8358)));
	track_2_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8361 downto 8360)));
	track_2_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8363 downto 8362)));
	track_2_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8365 downto 8364)));
	track_2_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8367 downto 8366)));
	track_2_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8369 downto 8368)));
	track_2_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8371 downto 8370)));
	track_2_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8373 downto 8372)));
	track_2_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8375 downto 8374)));
	track_2_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8377 downto 8376)));
	track_2_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8379 downto 8378)));
	track_2_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8381 downto 8380)));
	track_2_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8383 downto 8382)));
	track_2_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8385 downto 8384)));
	track_2_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8387 downto 8386)));
	track_2_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8389 downto 8388)));
	track_2_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8391 downto 8390)));
	track_2_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8393 downto 8392)));
	track_2_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8395 downto 8394)));
	track_2_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8397 downto 8396)));
	track_2_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8399 downto 8398)));
	track_2_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8401 downto 8400)));
	track_2_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8403 downto 8402)));
	track_2_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8405 downto 8404)));
	track_2_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8407 downto 8406)));
	track_2_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8409 downto 8408)));
	track_2_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8411 downto 8410)));
	track_2_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8413 downto 8412)));
	track_2_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8415 downto 8414)));
	track_2_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8417 downto 8416)));
	track_2_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8419 downto 8418)));
	track_2_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8421 downto 8420)));
	track_2_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8423 downto 8422)));
	track_2_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8425 downto 8424)));
	track_2_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8427 downto 8426)));
	track_2_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8429 downto 8428)));
	track_2_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8431 downto 8430)));
	track_2_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8433 downto 8432)));
	track_2_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8435 downto 8434)));
	track_2_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8437 downto 8436)));
	track_2_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8439 downto 8438)));
	track_2_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8441 downto 8440)));
	track_2_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8443 downto 8442)));
	track_2_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8445 downto 8444)));
	track_2_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8447 downto 8446)));
	track_2_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8449 downto 8448)));
	track_2_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8451 downto 8450)));
	track_2_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8453 downto 8452)));
	track_2_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8455 downto 8454)));
	track_2_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8457 downto 8456)));
	track_2_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8459 downto 8458)));
	track_2_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8461 downto 8460)));
	track_2_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8463 downto 8462)));
	track_2_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8465 downto 8464)));
	track_2_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8467 downto 8466)));
	track_2_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8469 downto 8468)));
	track_2_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8471 downto 8470)));
	track_3_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8473 downto 8472)));
	track_3_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8475 downto 8474)));
	track_3_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8477 downto 8476)));
	track_3_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8479 downto 8478)));
	track_3_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8481 downto 8480)));
	track_3_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8483 downto 8482)));
	track_3_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8485 downto 8484)));
	track_3_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8487 downto 8486)));
	track_3_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8489 downto 8488)));
	track_3_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8491 downto 8490)));
	track_3_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8493 downto 8492)));
	track_3_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8495 downto 8494)));
	track_3_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8497 downto 8496)));
	track_3_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8499 downto 8498)));
	track_3_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8501 downto 8500)));
	track_3_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8503 downto 8502)));
	track_3_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8505 downto 8504)));
	track_3_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8507 downto 8506)));
	track_3_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8509 downto 8508)));
	track_3_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8511 downto 8510)));
	track_3_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8513 downto 8512)));
	track_3_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8515 downto 8514)));
	track_3_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8517 downto 8516)));
	track_3_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8519 downto 8518)));
	track_3_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8521 downto 8520)));
	track_3_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8523 downto 8522)));
	track_3_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8525 downto 8524)));
	track_3_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8527 downto 8526)));
	track_3_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8529 downto 8528)));
	track_3_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8531 downto 8530)));
	track_3_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8533 downto 8532)));
	track_3_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8535 downto 8534)));
	track_3_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8537 downto 8536)));
	track_3_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8539 downto 8538)));
	track_3_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8541 downto 8540)));
	track_3_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8543 downto 8542)));
	track_3_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8545 downto 8544)));
	track_3_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8547 downto 8546)));
	track_3_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8549 downto 8548)));
	track_3_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8551 downto 8550)));
	track_3_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8553 downto 8552)));
	track_3_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8555 downto 8554)));
	track_3_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8557 downto 8556)));
	track_3_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8559 downto 8558)));
	track_3_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8561 downto 8560)));
	track_3_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8563 downto 8562)));
	track_3_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8565 downto 8564)));
	track_3_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8567 downto 8566)));
	track_3_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8569 downto 8568)));
	track_3_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8571 downto 8570)));
	track_3_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8573 downto 8572)));
	track_3_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8575 downto 8574)));
	track_3_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8577 downto 8576)));
	track_3_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8579 downto 8578)));
	track_3_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8581 downto 8580)));
	track_3_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8583 downto 8582)));
	track_3_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8585 downto 8584)));
	track_3_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8587 downto 8586)));
	track_3_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8589 downto 8588)));
	track_3_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8591 downto 8590)));
	track_3_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8593 downto 8592)));
	track_3_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8595 downto 8594)));
	track_3_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8597 downto 8596)));
	track_3_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8599 downto 8598)));
	track_3_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8601 downto 8600)));
	track_3_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8603 downto 8602)));
	track_3_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8605 downto 8604)));
	track_3_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8607 downto 8606)));
	track_3_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8609 downto 8608)));
	track_3_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8611 downto 8610)));
	track_3_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8613 downto 8612)));
	track_3_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8615 downto 8614)));
	track_3_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8617 downto 8616)));
	track_3_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8619 downto 8618)));
	track_3_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8621 downto 8620)));
	track_3_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8623 downto 8622)));
	track_3_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8625 downto 8624)));
	track_3_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8627 downto 8626)));
	track_3_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8629 downto 8628)));
	track_3_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8631 downto 8630)));
	track_3_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8633 downto 8632)));
	track_3_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8635 downto 8634)));
	track_3_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8637 downto 8636)));
	track_3_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8639 downto 8638)));
	track_3_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8641 downto 8640)));
	track_3_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8643 downto 8642)));
	track_3_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8645 downto 8644)));
	track_3_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8647 downto 8646)));
	track_3_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8649 downto 8648)));
	track_3_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8651 downto 8650)));
	track_3_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8653 downto 8652)));
	track_3_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8655 downto 8654)));
	track_3_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8657 downto 8656)));
	track_3_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8659 downto 8658)));
	track_3_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8661 downto 8660)));
	track_3_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8663 downto 8662)));
	track_3_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8665 downto 8664)));
	track_3_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8667 downto 8666)));
	track_3_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8669 downto 8668)));
	track_3_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8671 downto 8670)));
	track_3_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8673 downto 8672)));
	track_3_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8675 downto 8674)));
	track_3_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8677 downto 8676)));
	track_3_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8679 downto 8678)));
	track_3_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8681 downto 8680)));
	track_3_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8683 downto 8682)));
	track_3_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8685 downto 8684)));
	track_3_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8687 downto 8686)));
	track_3_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8689 downto 8688)));
	track_3_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8691 downto 8690)));
	track_3_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8693 downto 8692)));
	track_3_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8695 downto 8694)));
	track_3_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8697 downto 8696)));
	track_3_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8699 downto 8698)));
	track_3_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8701 downto 8700)));
	track_3_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8703 downto 8702)));
	track_3_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8705 downto 8704)));
	track_3_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8707 downto 8706)));
	track_3_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8709 downto 8708)));
	track_3_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8711 downto 8710)));
	track_3_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8713 downto 8712)));
	track_3_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8715 downto 8714)));
	track_3_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8717 downto 8716)));
	track_3_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8719 downto 8718)));
	track_3_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8721 downto 8720)));
	track_3_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8723 downto 8722)));
	track_3_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8725 downto 8724)));
	track_3_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8727 downto 8726)));
	track_3_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8729 downto 8728)));
	track_3_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8731 downto 8730)));
	track_3_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8733 downto 8732)));
	track_3_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8735 downto 8734)));
	track_3_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8737 downto 8736)));
	track_3_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8739 downto 8738)));
	track_3_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8741 downto 8740)));
	track_3_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8743 downto 8742)));
	track_3_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8745 downto 8744)));
	track_3_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8747 downto 8746)));
	track_3_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8749 downto 8748)));
	track_3_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8751 downto 8750)));
	track_3_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8753 downto 8752)));
	track_3_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8755 downto 8754)));
	track_3_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8757 downto 8756)));
	track_3_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8759 downto 8758)));
	track_3_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8761 downto 8760)));
	track_3_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8763 downto 8762)));
	track_3_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8765 downto 8764)));
	track_3_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8767 downto 8766)));
	track_3_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8769 downto 8768)));
	track_3_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8771 downto 8770)));
	track_3_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8773 downto 8772)));
	track_3_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8775 downto 8774)));
	track_3_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8777 downto 8776)));
	track_3_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8779 downto 8778)));
	track_3_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8781 downto 8780)));
	track_3_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8783 downto 8782)));
	track_3_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8785 downto 8784)));
	track_3_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8787 downto 8786)));
	track_3_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8789 downto 8788)));
	track_3_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8791 downto 8790)));
	track_3_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8793 downto 8792)));
	track_3_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8795 downto 8794)));
	track_3_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8797 downto 8796)));
	track_3_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8799 downto 8798)));
	track_3_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8801 downto 8800)));
	track_3_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8803 downto 8802)));
	track_3_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8805 downto 8804)));
	track_3_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8807 downto 8806)));
	track_3_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8809 downto 8808)));
	track_3_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8811 downto 8810)));
	track_3_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8813 downto 8812)));
	track_3_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8815 downto 8814)));
	track_3_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8817 downto 8816)));
	track_3_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8819 downto 8818)));
	track_3_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8821 downto 8820)));
	track_3_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8823 downto 8822)));
	track_3_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8825 downto 8824)));
	track_3_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8827 downto 8826)));
	track_3_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8829 downto 8828)));
	track_3_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8831 downto 8830)));
	track_3_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8833 downto 8832)));
	track_3_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8835 downto 8834)));
	track_3_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8837 downto 8836)));
	track_3_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8839 downto 8838)));
	track_3_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8841 downto 8840)));
	track_3_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8843 downto 8842)));
	track_3_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8845 downto 8844)));
	track_3_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8847 downto 8846)));
	track_3_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8849 downto 8848)));
	track_3_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8851 downto 8850)));
	track_3_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8853 downto 8852)));
	track_3_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8855 downto 8854)));
	track_3_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8857 downto 8856)));
	track_3_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8859 downto 8858)));
	track_3_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8861 downto 8860)));
	track_3_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8863 downto 8862)));
	track_3_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8865 downto 8864)));
	track_3_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8867 downto 8866)));
	track_3_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8869 downto 8868)));
	track_3_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8871 downto 8870)));
	track_3_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8873 downto 8872)));
	track_3_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8875 downto 8874)));
	track_3_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8877 downto 8876)));
	track_3_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8879 downto 8878)));
	track_3_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8881 downto 8880)));
	track_3_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8883 downto 8882)));
	track_3_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8885 downto 8884)));
	track_3_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8887 downto 8886)));
	track_4_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8889 downto 8888)));
	track_4_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8891 downto 8890)));
	track_4_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8893 downto 8892)));
	track_4_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8895 downto 8894)));
	track_4_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8897 downto 8896)));
	track_4_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8899 downto 8898)));
	track_4_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8901 downto 8900)));
	track_4_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8903 downto 8902)));
	track_4_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8905 downto 8904)));
	track_4_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8907 downto 8906)));
	track_4_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8909 downto 8908)));
	track_4_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8911 downto 8910)));
	track_4_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8913 downto 8912)));
	track_4_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8915 downto 8914)));
	track_4_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8917 downto 8916)));
	track_4_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8919 downto 8918)));
	track_4_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8921 downto 8920)));
	track_4_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8923 downto 8922)));
	track_4_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8925 downto 8924)));
	track_4_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8927 downto 8926)));
	track_4_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8929 downto 8928)));
	track_4_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8931 downto 8930)));
	track_4_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8933 downto 8932)));
	track_4_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8935 downto 8934)));
	track_4_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(8937 downto 8936)));
	track_4_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(8939 downto 8938)));
	track_4_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(8941 downto 8940)));
	track_4_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(8943 downto 8942)));
	track_4_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(8945 downto 8944)));
	track_4_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(8947 downto 8946)));
	track_4_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(8949 downto 8948)));
	track_4_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(8951 downto 8950)));
	track_4_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(8953 downto 8952)));
	track_4_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(8955 downto 8954)));
	track_4_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(8957 downto 8956)));
	track_4_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(8959 downto 8958)));
	track_4_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(8961 downto 8960)));
	track_4_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(8963 downto 8962)));
	track_4_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(8965 downto 8964)));
	track_4_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(8967 downto 8966)));
	track_4_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(8969 downto 8968)));
	track_4_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(8971 downto 8970)));
	track_4_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(8973 downto 8972)));
	track_4_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(8975 downto 8974)));
	track_4_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(8977 downto 8976)));
	track_4_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(8979 downto 8978)));
	track_4_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(8981 downto 8980)));
	track_4_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(8983 downto 8982)));
	track_4_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(8985 downto 8984)));
	track_4_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(8987 downto 8986)));
	track_4_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(8989 downto 8988)));
	track_4_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(8991 downto 8990)));
	track_4_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(8993 downto 8992)));
	track_4_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(8995 downto 8994)));
	track_4_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(8997 downto 8996)));
	track_4_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(8999 downto 8998)));
	track_4_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9001 downto 9000)));
	track_4_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9003 downto 9002)));
	track_4_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9005 downto 9004)));
	track_4_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9007 downto 9006)));
	track_4_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9009 downto 9008)));
	track_4_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9011 downto 9010)));
	track_4_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9013 downto 9012)));
	track_4_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9015 downto 9014)));
	track_4_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9017 downto 9016)));
	track_4_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9019 downto 9018)));
	track_4_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9021 downto 9020)));
	track_4_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9023 downto 9022)));
	track_4_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9025 downto 9024)));
	track_4_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9027 downto 9026)));
	track_4_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9029 downto 9028)));
	track_4_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9031 downto 9030)));
	track_4_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9033 downto 9032)));
	track_4_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9035 downto 9034)));
	track_4_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9037 downto 9036)));
	track_4_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9039 downto 9038)));
	track_4_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9041 downto 9040)));
	track_4_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9043 downto 9042)));
	track_4_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9045 downto 9044)));
	track_4_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9047 downto 9046)));
	track_4_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9049 downto 9048)));
	track_4_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9051 downto 9050)));
	track_4_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9053 downto 9052)));
	track_4_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9055 downto 9054)));
	track_4_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9057 downto 9056)));
	track_4_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9059 downto 9058)));
	track_4_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9061 downto 9060)));
	track_4_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9063 downto 9062)));
	track_4_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9065 downto 9064)));
	track_4_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9067 downto 9066)));
	track_4_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9069 downto 9068)));
	track_4_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9071 downto 9070)));
	track_4_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9073 downto 9072)));
	track_4_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9075 downto 9074)));
	track_4_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9077 downto 9076)));
	track_4_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9079 downto 9078)));
	track_4_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9081 downto 9080)));
	track_4_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9083 downto 9082)));
	track_4_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9085 downto 9084)));
	track_4_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9087 downto 9086)));
	track_4_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9089 downto 9088)));
	track_4_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9091 downto 9090)));
	track_4_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9093 downto 9092)));
	track_4_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9095 downto 9094)));
	track_4_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9097 downto 9096)));
	track_4_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9099 downto 9098)));
	track_4_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9101 downto 9100)));
	track_4_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9103 downto 9102)));
	track_4_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9105 downto 9104)));
	track_4_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9107 downto 9106)));
	track_4_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9109 downto 9108)));
	track_4_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9111 downto 9110)));
	track_4_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9113 downto 9112)));
	track_4_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9115 downto 9114)));
	track_4_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9117 downto 9116)));
	track_4_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9119 downto 9118)));
	track_4_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9121 downto 9120)));
	track_4_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9123 downto 9122)));
	track_4_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9125 downto 9124)));
	track_4_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9127 downto 9126)));
	track_4_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9129 downto 9128)));
	track_4_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9131 downto 9130)));
	track_4_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9133 downto 9132)));
	track_4_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9135 downto 9134)));
	track_4_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9137 downto 9136)));
	track_4_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9139 downto 9138)));
	track_4_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9141 downto 9140)));
	track_4_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9143 downto 9142)));
	track_4_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9145 downto 9144)));
	track_4_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9147 downto 9146)));
	track_4_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9149 downto 9148)));
	track_4_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9151 downto 9150)));
	track_4_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9153 downto 9152)));
	track_4_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9155 downto 9154)));
	track_4_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9157 downto 9156)));
	track_4_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9159 downto 9158)));
	track_4_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9161 downto 9160)));
	track_4_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9163 downto 9162)));
	track_4_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9165 downto 9164)));
	track_4_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9167 downto 9166)));
	track_4_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9169 downto 9168)));
	track_4_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9171 downto 9170)));
	track_4_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9173 downto 9172)));
	track_4_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9175 downto 9174)));
	track_4_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9177 downto 9176)));
	track_4_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9179 downto 9178)));
	track_4_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9181 downto 9180)));
	track_4_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9183 downto 9182)));
	track_4_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9185 downto 9184)));
	track_4_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9187 downto 9186)));
	track_4_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9189 downto 9188)));
	track_4_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9191 downto 9190)));
	track_4_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9193 downto 9192)));
	track_4_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9195 downto 9194)));
	track_4_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9197 downto 9196)));
	track_4_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9199 downto 9198)));
	track_4_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9201 downto 9200)));
	track_4_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9203 downto 9202)));
	track_4_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9205 downto 9204)));
	track_4_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9207 downto 9206)));
	track_4_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9209 downto 9208)));
	track_4_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9211 downto 9210)));
	track_4_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9213 downto 9212)));
	track_4_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9215 downto 9214)));
	track_4_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9217 downto 9216)));
	track_4_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9219 downto 9218)));
	track_4_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9221 downto 9220)));
	track_4_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9223 downto 9222)));
	track_4_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9225 downto 9224)));
	track_4_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9227 downto 9226)));
	track_4_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9229 downto 9228)));
	track_4_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9231 downto 9230)));
	track_4_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9233 downto 9232)));
	track_4_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9235 downto 9234)));
	track_4_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9237 downto 9236)));
	track_4_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9239 downto 9238)));
	track_4_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9241 downto 9240)));
	track_4_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9243 downto 9242)));
	track_4_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9245 downto 9244)));
	track_4_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9247 downto 9246)));
	track_4_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9249 downto 9248)));
	track_4_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9251 downto 9250)));
	track_4_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9253 downto 9252)));
	track_4_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9255 downto 9254)));
	track_4_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9257 downto 9256)));
	track_4_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9259 downto 9258)));
	track_4_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9261 downto 9260)));
	track_4_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9263 downto 9262)));
	track_4_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9265 downto 9264)));
	track_4_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9267 downto 9266)));
	track_4_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9269 downto 9268)));
	track_4_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9271 downto 9270)));
	track_4_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9273 downto 9272)));
	track_4_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9275 downto 9274)));
	track_4_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9277 downto 9276)));
	track_4_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9279 downto 9278)));
	track_4_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9281 downto 9280)));
	track_4_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9283 downto 9282)));
	track_4_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9285 downto 9284)));
	track_4_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9287 downto 9286)));
	track_4_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9289 downto 9288)));
	track_4_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9291 downto 9290)));
	track_4_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9293 downto 9292)));
	track_4_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9295 downto 9294)));
	track_4_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9297 downto 9296)));
	track_4_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9299 downto 9298)));
	track_4_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9301 downto 9300)));
	track_4_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9303 downto 9302)));
	track_5_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9305 downto 9304)));
	track_5_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9307 downto 9306)));
	track_5_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9309 downto 9308)));
	track_5_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9311 downto 9310)));
	track_5_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9313 downto 9312)));
	track_5_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9315 downto 9314)));
	track_5_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9317 downto 9316)));
	track_5_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9319 downto 9318)));
	track_5_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9321 downto 9320)));
	track_5_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9323 downto 9322)));
	track_5_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9325 downto 9324)));
	track_5_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9327 downto 9326)));
	track_5_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9329 downto 9328)));
	track_5_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9331 downto 9330)));
	track_5_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9333 downto 9332)));
	track_5_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9335 downto 9334)));
	track_5_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9337 downto 9336)));
	track_5_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9339 downto 9338)));
	track_5_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9341 downto 9340)));
	track_5_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9343 downto 9342)));
	track_5_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9345 downto 9344)));
	track_5_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9347 downto 9346)));
	track_5_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9349 downto 9348)));
	track_5_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9351 downto 9350)));
	track_5_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9353 downto 9352)));
	track_5_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9355 downto 9354)));
	track_5_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9357 downto 9356)));
	track_5_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9359 downto 9358)));
	track_5_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9361 downto 9360)));
	track_5_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9363 downto 9362)));
	track_5_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9365 downto 9364)));
	track_5_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9367 downto 9366)));
	track_5_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9369 downto 9368)));
	track_5_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9371 downto 9370)));
	track_5_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9373 downto 9372)));
	track_5_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9375 downto 9374)));
	track_5_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9377 downto 9376)));
	track_5_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9379 downto 9378)));
	track_5_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9381 downto 9380)));
	track_5_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9383 downto 9382)));
	track_5_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9385 downto 9384)));
	track_5_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9387 downto 9386)));
	track_5_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9389 downto 9388)));
	track_5_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9391 downto 9390)));
	track_5_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9393 downto 9392)));
	track_5_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9395 downto 9394)));
	track_5_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9397 downto 9396)));
	track_5_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9399 downto 9398)));
	track_5_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9401 downto 9400)));
	track_5_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9403 downto 9402)));
	track_5_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9405 downto 9404)));
	track_5_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9407 downto 9406)));
	track_5_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9409 downto 9408)));
	track_5_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9411 downto 9410)));
	track_5_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9413 downto 9412)));
	track_5_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9415 downto 9414)));
	track_5_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9417 downto 9416)));
	track_5_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9419 downto 9418)));
	track_5_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9421 downto 9420)));
	track_5_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9423 downto 9422)));
	track_5_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9425 downto 9424)));
	track_5_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9427 downto 9426)));
	track_5_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9429 downto 9428)));
	track_5_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9431 downto 9430)));
	track_5_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9433 downto 9432)));
	track_5_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9435 downto 9434)));
	track_5_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9437 downto 9436)));
	track_5_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9439 downto 9438)));
	track_5_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9441 downto 9440)));
	track_5_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9443 downto 9442)));
	track_5_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9445 downto 9444)));
	track_5_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9447 downto 9446)));
	track_5_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9449 downto 9448)));
	track_5_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9451 downto 9450)));
	track_5_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9453 downto 9452)));
	track_5_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9455 downto 9454)));
	track_5_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9457 downto 9456)));
	track_5_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9459 downto 9458)));
	track_5_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9461 downto 9460)));
	track_5_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9463 downto 9462)));
	track_5_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9465 downto 9464)));
	track_5_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9467 downto 9466)));
	track_5_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9469 downto 9468)));
	track_5_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9471 downto 9470)));
	track_5_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9473 downto 9472)));
	track_5_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9475 downto 9474)));
	track_5_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9477 downto 9476)));
	track_5_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9479 downto 9478)));
	track_5_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9481 downto 9480)));
	track_5_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9483 downto 9482)));
	track_5_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9485 downto 9484)));
	track_5_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9487 downto 9486)));
	track_5_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9489 downto 9488)));
	track_5_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9491 downto 9490)));
	track_5_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9493 downto 9492)));
	track_5_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9495 downto 9494)));
	track_5_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9497 downto 9496)));
	track_5_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9499 downto 9498)));
	track_5_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9501 downto 9500)));
	track_5_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9503 downto 9502)));
	track_5_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9505 downto 9504)));
	track_5_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9507 downto 9506)));
	track_5_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9509 downto 9508)));
	track_5_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9511 downto 9510)));
	track_5_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9513 downto 9512)));
	track_5_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9515 downto 9514)));
	track_5_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9517 downto 9516)));
	track_5_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9519 downto 9518)));
	track_5_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9521 downto 9520)));
	track_5_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9523 downto 9522)));
	track_5_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9525 downto 9524)));
	track_5_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9527 downto 9526)));
	track_5_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9529 downto 9528)));
	track_5_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9531 downto 9530)));
	track_5_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9533 downto 9532)));
	track_5_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9535 downto 9534)));
	track_5_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9537 downto 9536)));
	track_5_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9539 downto 9538)));
	track_5_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9541 downto 9540)));
	track_5_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9543 downto 9542)));
	track_5_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9545 downto 9544)));
	track_5_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9547 downto 9546)));
	track_5_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9549 downto 9548)));
	track_5_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9551 downto 9550)));
	track_5_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9553 downto 9552)));
	track_5_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9555 downto 9554)));
	track_5_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9557 downto 9556)));
	track_5_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9559 downto 9558)));
	track_5_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9561 downto 9560)));
	track_5_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9563 downto 9562)));
	track_5_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9565 downto 9564)));
	track_5_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9567 downto 9566)));
	track_5_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9569 downto 9568)));
	track_5_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9571 downto 9570)));
	track_5_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9573 downto 9572)));
	track_5_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9575 downto 9574)));
	track_5_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9577 downto 9576)));
	track_5_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9579 downto 9578)));
	track_5_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9581 downto 9580)));
	track_5_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9583 downto 9582)));
	track_5_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9585 downto 9584)));
	track_5_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9587 downto 9586)));
	track_5_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9589 downto 9588)));
	track_5_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9591 downto 9590)));
	track_5_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9593 downto 9592)));
	track_5_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9595 downto 9594)));
	track_5_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9597 downto 9596)));
	track_5_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9599 downto 9598)));
	track_5_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9601 downto 9600)));
	track_5_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9603 downto 9602)));
	track_5_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9605 downto 9604)));
	track_5_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9607 downto 9606)));
	track_5_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9609 downto 9608)));
	track_5_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9611 downto 9610)));
	track_5_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9613 downto 9612)));
	track_5_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9615 downto 9614)));
	track_5_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9617 downto 9616)));
	track_5_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9619 downto 9618)));
	track_5_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9621 downto 9620)));
	track_5_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9623 downto 9622)));
	track_5_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9625 downto 9624)));
	track_5_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9627 downto 9626)));
	track_5_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9629 downto 9628)));
	track_5_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9631 downto 9630)));
	track_5_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9633 downto 9632)));
	track_5_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9635 downto 9634)));
	track_5_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9637 downto 9636)));
	track_5_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9639 downto 9638)));
	track_5_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9641 downto 9640)));
	track_5_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9643 downto 9642)));
	track_5_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9645 downto 9644)));
	track_5_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9647 downto 9646)));
	track_5_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9649 downto 9648)));
	track_5_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9651 downto 9650)));
	track_5_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9653 downto 9652)));
	track_5_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9655 downto 9654)));
	track_5_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9657 downto 9656)));
	track_5_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9659 downto 9658)));
	track_5_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9661 downto 9660)));
	track_5_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9663 downto 9662)));
	track_5_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9665 downto 9664)));
	track_5_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9667 downto 9666)));
	track_5_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9669 downto 9668)));
	track_5_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9671 downto 9670)));
	track_5_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9673 downto 9672)));
	track_5_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9675 downto 9674)));
	track_5_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9677 downto 9676)));
	track_5_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9679 downto 9678)));
	track_5_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9681 downto 9680)));
	track_5_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9683 downto 9682)));
	track_5_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9685 downto 9684)));
	track_5_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9687 downto 9686)));
	track_5_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9689 downto 9688)));
	track_5_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9691 downto 9690)));
	track_5_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9693 downto 9692)));
	track_5_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9695 downto 9694)));
	track_5_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9697 downto 9696)));
	track_5_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9699 downto 9698)));
	track_5_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9701 downto 9700)));
	track_5_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9703 downto 9702)));
	track_5_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9705 downto 9704)));
	track_5_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9707 downto 9706)));
	track_5_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9709 downto 9708)));
	track_5_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9711 downto 9710)));
	track_5_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9713 downto 9712)));
	track_5_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9715 downto 9714)));
	track_5_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9717 downto 9716)));
	track_5_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9719 downto 9718)));
	track_6_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9721 downto 9720)));
	track_6_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9723 downto 9722)));
	track_6_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9725 downto 9724)));
	track_6_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9727 downto 9726)));
	track_6_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9729 downto 9728)));
	track_6_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9731 downto 9730)));
	track_6_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9733 downto 9732)));
	track_6_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9735 downto 9734)));
	track_6_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9737 downto 9736)));
	track_6_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9739 downto 9738)));
	track_6_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9741 downto 9740)));
	track_6_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9743 downto 9742)));
	track_6_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9745 downto 9744)));
	track_6_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9747 downto 9746)));
	track_6_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9749 downto 9748)));
	track_6_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9751 downto 9750)));
	track_6_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9753 downto 9752)));
	track_6_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9755 downto 9754)));
	track_6_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9757 downto 9756)));
	track_6_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9759 downto 9758)));
	track_6_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9761 downto 9760)));
	track_6_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9763 downto 9762)));
	track_6_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9765 downto 9764)));
	track_6_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9767 downto 9766)));
	track_6_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9769 downto 9768)));
	track_6_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9771 downto 9770)));
	track_6_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9773 downto 9772)));
	track_6_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9775 downto 9774)));
	track_6_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9777 downto 9776)));
	track_6_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9779 downto 9778)));
	track_6_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9781 downto 9780)));
	track_6_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9783 downto 9782)));
	track_6_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9785 downto 9784)));
	track_6_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9787 downto 9786)));
	track_6_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9789 downto 9788)));
	track_6_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9791 downto 9790)));
	track_6_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9793 downto 9792)));
	track_6_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9795 downto 9794)));
	track_6_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9797 downto 9796)));
	track_6_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9799 downto 9798)));
	track_6_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9801 downto 9800)));
	track_6_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9803 downto 9802)));
	track_6_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9805 downto 9804)));
	track_6_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9807 downto 9806)));
	track_6_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9809 downto 9808)));
	track_6_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9811 downto 9810)));
	track_6_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9813 downto 9812)));
	track_6_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9815 downto 9814)));
	track_6_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9817 downto 9816)));
	track_6_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9819 downto 9818)));
	track_6_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9821 downto 9820)));
	track_6_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9823 downto 9822)));
	track_6_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9825 downto 9824)));
	track_6_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9827 downto 9826)));
	track_6_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9829 downto 9828)));
	track_6_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9831 downto 9830)));
	track_6_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9833 downto 9832)));
	track_6_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9835 downto 9834)));
	track_6_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9837 downto 9836)));
	track_6_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9839 downto 9838)));
	track_6_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9841 downto 9840)));
	track_6_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9843 downto 9842)));
	track_6_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9845 downto 9844)));
	track_6_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9847 downto 9846)));
	track_6_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9849 downto 9848)));
	track_6_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9851 downto 9850)));
	track_6_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9853 downto 9852)));
	track_6_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9855 downto 9854)));
	track_6_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9857 downto 9856)));
	track_6_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9859 downto 9858)));
	track_6_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9861 downto 9860)));
	track_6_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9863 downto 9862)));
	track_6_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9865 downto 9864)));
	track_6_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9867 downto 9866)));
	track_6_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9869 downto 9868)));
	track_6_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9871 downto 9870)));
	track_6_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9873 downto 9872)));
	track_6_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9875 downto 9874)));
	track_6_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9877 downto 9876)));
	track_6_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9879 downto 9878)));
	track_6_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9881 downto 9880)));
	track_6_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9883 downto 9882)));
	track_6_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9885 downto 9884)));
	track_6_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9887 downto 9886)));
	track_6_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9889 downto 9888)));
	track_6_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9891 downto 9890)));
	track_6_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9893 downto 9892)));
	track_6_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9895 downto 9894)));
	track_6_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9897 downto 9896)));
	track_6_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9899 downto 9898)));
	track_6_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9901 downto 9900)));
	track_6_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9903 downto 9902)));
	track_6_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9905 downto 9904)));
	track_6_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9907 downto 9906)));
	track_6_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9909 downto 9908)));
	track_6_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9911 downto 9910)));
	track_6_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9913 downto 9912)));
	track_6_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9915 downto 9914)));
	track_6_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9917 downto 9916)));
	track_6_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9919 downto 9918)));
	track_6_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9921 downto 9920)));
	track_6_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9923 downto 9922)));
	track_6_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9925 downto 9924)));
	track_6_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9927 downto 9926)));
	track_6_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9929 downto 9928)));
	track_6_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9931 downto 9930)));
	track_6_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9933 downto 9932)));
	track_6_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9935 downto 9934)));
	track_6_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(9937 downto 9936)));
	track_6_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(9939 downto 9938)));
	track_6_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(9941 downto 9940)));
	track_6_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(9943 downto 9942)));
	track_6_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(9945 downto 9944)));
	track_6_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(9947 downto 9946)));
	track_6_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(9949 downto 9948)));
	track_6_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(9951 downto 9950)));
	track_6_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(9953 downto 9952)));
	track_6_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(9955 downto 9954)));
	track_6_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(9957 downto 9956)));
	track_6_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(9959 downto 9958)));
	track_6_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(9961 downto 9960)));
	track_6_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(9963 downto 9962)));
	track_6_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(9965 downto 9964)));
	track_6_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(9967 downto 9966)));
	track_6_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(9969 downto 9968)));
	track_6_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(9971 downto 9970)));
	track_6_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(9973 downto 9972)));
	track_6_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(9975 downto 9974)));
	track_6_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(9977 downto 9976)));
	track_6_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(9979 downto 9978)));
	track_6_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(9981 downto 9980)));
	track_6_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(9983 downto 9982)));
	track_6_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(9985 downto 9984)));
	track_6_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(9987 downto 9986)));
	track_6_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(9989 downto 9988)));
	track_6_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(9991 downto 9990)));
	track_6_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(9993 downto 9992)));
	track_6_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(9995 downto 9994)));
	track_6_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(9997 downto 9996)));
	track_6_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(9999 downto 9998)));
	track_6_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10001 downto 10000)));
	track_6_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10003 downto 10002)));
	track_6_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10005 downto 10004)));
	track_6_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10007 downto 10006)));
	track_6_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10009 downto 10008)));
	track_6_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10011 downto 10010)));
	track_6_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10013 downto 10012)));
	track_6_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10015 downto 10014)));
	track_6_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10017 downto 10016)));
	track_6_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10019 downto 10018)));
	track_6_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10021 downto 10020)));
	track_6_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10023 downto 10022)));
	track_6_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10025 downto 10024)));
	track_6_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10027 downto 10026)));
	track_6_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10029 downto 10028)));
	track_6_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10031 downto 10030)));
	track_6_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10033 downto 10032)));
	track_6_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10035 downto 10034)));
	track_6_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10037 downto 10036)));
	track_6_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10039 downto 10038)));
	track_6_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10041 downto 10040)));
	track_6_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10043 downto 10042)));
	track_6_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10045 downto 10044)));
	track_6_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10047 downto 10046)));
	track_6_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10049 downto 10048)));
	track_6_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10051 downto 10050)));
	track_6_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10053 downto 10052)));
	track_6_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10055 downto 10054)));
	track_6_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10057 downto 10056)));
	track_6_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10059 downto 10058)));
	track_6_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10061 downto 10060)));
	track_6_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10063 downto 10062)));
	track_6_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10065 downto 10064)));
	track_6_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10067 downto 10066)));
	track_6_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10069 downto 10068)));
	track_6_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10071 downto 10070)));
	track_6_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10073 downto 10072)));
	track_6_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10075 downto 10074)));
	track_6_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10077 downto 10076)));
	track_6_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10079 downto 10078)));
	track_6_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10081 downto 10080)));
	track_6_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10083 downto 10082)));
	track_6_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10085 downto 10084)));
	track_6_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10087 downto 10086)));
	track_6_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10089 downto 10088)));
	track_6_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10091 downto 10090)));
	track_6_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10093 downto 10092)));
	track_6_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10095 downto 10094)));
	track_6_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10097 downto 10096)));
	track_6_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10099 downto 10098)));
	track_6_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10101 downto 10100)));
	track_6_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10103 downto 10102)));
	track_6_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10105 downto 10104)));
	track_6_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10107 downto 10106)));
	track_6_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10109 downto 10108)));
	track_6_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10111 downto 10110)));
	track_6_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10113 downto 10112)));
	track_6_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10115 downto 10114)));
	track_6_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10117 downto 10116)));
	track_6_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10119 downto 10118)));
	track_6_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10121 downto 10120)));
	track_6_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10123 downto 10122)));
	track_6_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10125 downto 10124)));
	track_6_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10127 downto 10126)));
	track_6_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10129 downto 10128)));
	track_6_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10131 downto 10130)));
	track_6_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10133 downto 10132)));
	track_6_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10135 downto 10134)));
	track_7_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10137 downto 10136)));
	track_7_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10139 downto 10138)));
	track_7_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10141 downto 10140)));
	track_7_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10143 downto 10142)));
	track_7_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10145 downto 10144)));
	track_7_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10147 downto 10146)));
	track_7_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10149 downto 10148)));
	track_7_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10151 downto 10150)));
	track_7_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10153 downto 10152)));
	track_7_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10155 downto 10154)));
	track_7_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10157 downto 10156)));
	track_7_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10159 downto 10158)));
	track_7_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10161 downto 10160)));
	track_7_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10163 downto 10162)));
	track_7_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10165 downto 10164)));
	track_7_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10167 downto 10166)));
	track_7_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10169 downto 10168)));
	track_7_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10171 downto 10170)));
	track_7_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10173 downto 10172)));
	track_7_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10175 downto 10174)));
	track_7_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10177 downto 10176)));
	track_7_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10179 downto 10178)));
	track_7_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10181 downto 10180)));
	track_7_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10183 downto 10182)));
	track_7_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10185 downto 10184)));
	track_7_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10187 downto 10186)));
	track_7_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10189 downto 10188)));
	track_7_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10191 downto 10190)));
	track_7_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10193 downto 10192)));
	track_7_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10195 downto 10194)));
	track_7_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10197 downto 10196)));
	track_7_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10199 downto 10198)));
	track_7_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10201 downto 10200)));
	track_7_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10203 downto 10202)));
	track_7_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10205 downto 10204)));
	track_7_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10207 downto 10206)));
	track_7_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10209 downto 10208)));
	track_7_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10211 downto 10210)));
	track_7_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10213 downto 10212)));
	track_7_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10215 downto 10214)));
	track_7_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10217 downto 10216)));
	track_7_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10219 downto 10218)));
	track_7_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10221 downto 10220)));
	track_7_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10223 downto 10222)));
	track_7_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10225 downto 10224)));
	track_7_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10227 downto 10226)));
	track_7_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10229 downto 10228)));
	track_7_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10231 downto 10230)));
	track_7_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10233 downto 10232)));
	track_7_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10235 downto 10234)));
	track_7_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10237 downto 10236)));
	track_7_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10239 downto 10238)));
	track_7_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10241 downto 10240)));
	track_7_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10243 downto 10242)));
	track_7_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10245 downto 10244)));
	track_7_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10247 downto 10246)));
	track_7_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10249 downto 10248)));
	track_7_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10251 downto 10250)));
	track_7_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10253 downto 10252)));
	track_7_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10255 downto 10254)));
	track_7_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10257 downto 10256)));
	track_7_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10259 downto 10258)));
	track_7_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10261 downto 10260)));
	track_7_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10263 downto 10262)));
	track_7_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10265 downto 10264)));
	track_7_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10267 downto 10266)));
	track_7_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10269 downto 10268)));
	track_7_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10271 downto 10270)));
	track_7_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10273 downto 10272)));
	track_7_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10275 downto 10274)));
	track_7_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10277 downto 10276)));
	track_7_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10279 downto 10278)));
	track_7_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10281 downto 10280)));
	track_7_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10283 downto 10282)));
	track_7_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10285 downto 10284)));
	track_7_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10287 downto 10286)));
	track_7_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10289 downto 10288)));
	track_7_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10291 downto 10290)));
	track_7_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10293 downto 10292)));
	track_7_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10295 downto 10294)));
	track_7_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10297 downto 10296)));
	track_7_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10299 downto 10298)));
	track_7_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10301 downto 10300)));
	track_7_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10303 downto 10302)));
	track_7_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10305 downto 10304)));
	track_7_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10307 downto 10306)));
	track_7_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10309 downto 10308)));
	track_7_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10311 downto 10310)));
	track_7_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10313 downto 10312)));
	track_7_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10315 downto 10314)));
	track_7_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10317 downto 10316)));
	track_7_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10319 downto 10318)));
	track_7_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10321 downto 10320)));
	track_7_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10323 downto 10322)));
	track_7_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10325 downto 10324)));
	track_7_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10327 downto 10326)));
	track_7_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10329 downto 10328)));
	track_7_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10331 downto 10330)));
	track_7_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10333 downto 10332)));
	track_7_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10335 downto 10334)));
	track_7_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10337 downto 10336)));
	track_7_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10339 downto 10338)));
	track_7_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10341 downto 10340)));
	track_7_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10343 downto 10342)));
	track_7_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10345 downto 10344)));
	track_7_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10347 downto 10346)));
	track_7_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10349 downto 10348)));
	track_7_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10351 downto 10350)));
	track_7_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10353 downto 10352)));
	track_7_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10355 downto 10354)));
	track_7_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10357 downto 10356)));
	track_7_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10359 downto 10358)));
	track_7_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10361 downto 10360)));
	track_7_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10363 downto 10362)));
	track_7_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10365 downto 10364)));
	track_7_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10367 downto 10366)));
	track_7_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10369 downto 10368)));
	track_7_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10371 downto 10370)));
	track_7_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10373 downto 10372)));
	track_7_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10375 downto 10374)));
	track_7_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10377 downto 10376)));
	track_7_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10379 downto 10378)));
	track_7_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10381 downto 10380)));
	track_7_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10383 downto 10382)));
	track_7_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10385 downto 10384)));
	track_7_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10387 downto 10386)));
	track_7_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10389 downto 10388)));
	track_7_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10391 downto 10390)));
	track_7_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10393 downto 10392)));
	track_7_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10395 downto 10394)));
	track_7_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10397 downto 10396)));
	track_7_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10399 downto 10398)));
	track_7_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10401 downto 10400)));
	track_7_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10403 downto 10402)));
	track_7_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10405 downto 10404)));
	track_7_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10407 downto 10406)));
	track_7_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10409 downto 10408)));
	track_7_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10411 downto 10410)));
	track_7_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10413 downto 10412)));
	track_7_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10415 downto 10414)));
	track_7_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10417 downto 10416)));
	track_7_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10419 downto 10418)));
	track_7_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10421 downto 10420)));
	track_7_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10423 downto 10422)));
	track_7_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10425 downto 10424)));
	track_7_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10427 downto 10426)));
	track_7_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10429 downto 10428)));
	track_7_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10431 downto 10430)));
	track_7_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10433 downto 10432)));
	track_7_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10435 downto 10434)));
	track_7_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10437 downto 10436)));
	track_7_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10439 downto 10438)));
	track_7_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10441 downto 10440)));
	track_7_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10443 downto 10442)));
	track_7_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10445 downto 10444)));
	track_7_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10447 downto 10446)));
	track_7_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10449 downto 10448)));
	track_7_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10451 downto 10450)));
	track_7_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10453 downto 10452)));
	track_7_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10455 downto 10454)));
	track_7_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10457 downto 10456)));
	track_7_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10459 downto 10458)));
	track_7_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10461 downto 10460)));
	track_7_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10463 downto 10462)));
	track_7_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10465 downto 10464)));
	track_7_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10467 downto 10466)));
	track_7_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10469 downto 10468)));
	track_7_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10471 downto 10470)));
	track_7_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10473 downto 10472)));
	track_7_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10475 downto 10474)));
	track_7_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10477 downto 10476)));
	track_7_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10479 downto 10478)));
	track_7_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10481 downto 10480)));
	track_7_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10483 downto 10482)));
	track_7_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10485 downto 10484)));
	track_7_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10487 downto 10486)));
	track_7_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10489 downto 10488)));
	track_7_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10491 downto 10490)));
	track_7_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10493 downto 10492)));
	track_7_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10495 downto 10494)));
	track_7_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10497 downto 10496)));
	track_7_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10499 downto 10498)));
	track_7_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10501 downto 10500)));
	track_7_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10503 downto 10502)));
	track_7_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10505 downto 10504)));
	track_7_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10507 downto 10506)));
	track_7_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10509 downto 10508)));
	track_7_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10511 downto 10510)));
	track_7_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10513 downto 10512)));
	track_7_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10515 downto 10514)));
	track_7_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10517 downto 10516)));
	track_7_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10519 downto 10518)));
	track_7_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10521 downto 10520)));
	track_7_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10523 downto 10522)));
	track_7_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10525 downto 10524)));
	track_7_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10527 downto 10526)));
	track_7_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10529 downto 10528)));
	track_7_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10531 downto 10530)));
	track_7_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10533 downto 10532)));
	track_7_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10535 downto 10534)));
	track_7_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10537 downto 10536)));
	track_7_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10539 downto 10538)));
	track_7_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10541 downto 10540)));
	track_7_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10543 downto 10542)));
	track_7_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10545 downto 10544)));
	track_7_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10547 downto 10546)));
	track_7_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10549 downto 10548)));
	track_7_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10551 downto 10550)));
	track_8_0_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10553 downto 10552)));
	track_8_0_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10555 downto 10554)));
	track_8_0_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10557 downto 10556)));
	track_8_0_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10558 downto 10558)));
	track_8_0_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10560 downto 10559)));
	track_8_0_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10561 downto 10561)));
	track_8_0_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10563 downto 10562)));
	track_8_0_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10564 downto 10564)));
	track_8_0_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10566 downto 10565)));
	track_8_0_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10568 downto 10567)));
	track_8_0_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10570 downto 10569)));
	track_8_0_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10572 downto 10571)));
	track_8_0_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10574 downto 10573)));
	track_8_0_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10576 downto 10575)));
	track_8_0_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10578 downto 10577)));
	track_8_0_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10579 downto 10579)));
	track_8_1_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10581 downto 10580)));
	track_8_1_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10583 downto 10582)));
	track_8_1_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10585 downto 10584)));
	track_8_1_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10587 downto 10586)));
	track_8_1_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10589 downto 10588)));
	track_8_1_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10591 downto 10590)));
	track_8_1_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10593 downto 10592)));
	track_8_1_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10595 downto 10594)));
	track_8_1_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10597 downto 10596)));
	track_8_1_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10599 downto 10598)));
	track_8_1_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10601 downto 10600)));
	track_8_1_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10603 downto 10602)));
	track_8_1_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10605 downto 10604)));
	track_8_1_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10607 downto 10606)));
	track_8_1_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10609 downto 10608)));
	track_8_1_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10611 downto 10610)));
	track_8_1_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10613 downto 10612)));
	track_8_1_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10615 downto 10614)));
	track_8_1_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10616 downto 10616)));
	track_8_1_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10618 downto 10617)));
	track_8_1_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10619 downto 10619)));
	track_8_1_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10621 downto 10620)));
	track_8_1_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10622 downto 10622)));
	track_8_1_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10624 downto 10623)));
	track_8_1_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10626 downto 10625)));
	track_8_1_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10628 downto 10627)));
	track_8_1_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10630 downto 10629)));
	track_8_1_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10632 downto 10631)));
	track_8_1_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10634 downto 10633)));
	track_8_1_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10636 downto 10635)));
	track_8_1_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10637 downto 10637)));
	track_8_1_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10639 downto 10638)));
	track_8_2_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10641 downto 10640)));
	track_8_2_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10643 downto 10642)));
	track_8_2_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10645 downto 10644)));
	track_8_2_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10647 downto 10646)));
	track_8_2_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10649 downto 10648)));
	track_8_2_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10651 downto 10650)));
	track_8_2_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10653 downto 10652)));
	track_8_2_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10655 downto 10654)));
	track_8_2_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10657 downto 10656)));
	track_8_2_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10659 downto 10658)));
	track_8_2_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10661 downto 10660)));
	track_8_2_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10663 downto 10662)));
	track_8_2_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10665 downto 10664)));
	track_8_2_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10667 downto 10666)));
	track_8_2_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10669 downto 10668)));
	track_8_2_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10671 downto 10670)));
	track_8_2_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10673 downto 10672)));
	track_8_2_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10675 downto 10674)));
	track_8_2_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10677 downto 10676)));
	track_8_2_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10679 downto 10678)));
	track_8_2_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10681 downto 10680)));
	track_8_2_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10683 downto 10682)));
	track_8_2_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10685 downto 10684)));
	track_8_2_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10687 downto 10686)));
	track_8_2_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10689 downto 10688)));
	track_8_2_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10691 downto 10690)));
	track_8_2_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10693 downto 10692)));
	track_8_2_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10695 downto 10694)));
	track_8_2_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10697 downto 10696)));
	track_8_2_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10699 downto 10698)));
	track_8_2_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10701 downto 10700)));
	track_8_2_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10703 downto 10702)));
	track_8_3_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10705 downto 10704)));
	track_8_3_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10707 downto 10706)));
	track_8_3_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10709 downto 10708)));
	track_8_3_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10711 downto 10710)));
	track_8_3_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10713 downto 10712)));
	track_8_3_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10715 downto 10714)));
	track_8_3_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10717 downto 10716)));
	track_8_3_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10719 downto 10718)));
	track_8_3_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10721 downto 10720)));
	track_8_3_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10723 downto 10722)));
	track_8_3_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10725 downto 10724)));
	track_8_3_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10727 downto 10726)));
	track_8_3_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10729 downto 10728)));
	track_8_3_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10731 downto 10730)));
	track_8_3_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10733 downto 10732)));
	track_8_3_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10735 downto 10734)));
	track_8_3_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10737 downto 10736)));
	track_8_3_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10739 downto 10738)));
	track_8_3_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10741 downto 10740)));
	track_8_3_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10743 downto 10742)));
	track_8_3_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10745 downto 10744)));
	track_8_3_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10747 downto 10746)));
	track_8_3_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10749 downto 10748)));
	track_8_3_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10751 downto 10750)));
	track_8_3_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10753 downto 10752)));
	track_8_3_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10755 downto 10754)));
	track_8_3_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10757 downto 10756)));
	track_8_3_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10759 downto 10758)));
	track_8_3_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10761 downto 10760)));
	track_8_3_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10763 downto 10762)));
	track_8_3_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10765 downto 10764)));
	track_8_3_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10767 downto 10766)));
	track_8_4_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10769 downto 10768)));
	track_8_4_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10771 downto 10770)));
	track_8_4_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10773 downto 10772)));
	track_8_4_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10775 downto 10774)));
	track_8_4_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10777 downto 10776)));
	track_8_4_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10779 downto 10778)));
	track_8_4_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10781 downto 10780)));
	track_8_4_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10783 downto 10782)));
	track_8_4_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10785 downto 10784)));
	track_8_4_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10787 downto 10786)));
	track_8_4_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10789 downto 10788)));
	track_8_4_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10791 downto 10790)));
	track_8_4_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10793 downto 10792)));
	track_8_4_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10795 downto 10794)));
	track_8_4_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10797 downto 10796)));
	track_8_4_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10799 downto 10798)));
	track_8_4_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10801 downto 10800)));
	track_8_4_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10803 downto 10802)));
	track_8_4_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10805 downto 10804)));
	track_8_4_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10807 downto 10806)));
	track_8_4_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10809 downto 10808)));
	track_8_4_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10811 downto 10810)));
	track_8_4_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10813 downto 10812)));
	track_8_4_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10815 downto 10814)));
	track_8_4_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10817 downto 10816)));
	track_8_4_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10819 downto 10818)));
	track_8_4_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10821 downto 10820)));
	track_8_4_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10823 downto 10822)));
	track_8_4_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10825 downto 10824)));
	track_8_4_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10827 downto 10826)));
	track_8_4_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10829 downto 10828)));
	track_8_4_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10831 downto 10830)));
	track_8_5_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10833 downto 10832)));
	track_8_5_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10835 downto 10834)));
	track_8_5_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10837 downto 10836)));
	track_8_5_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10839 downto 10838)));
	track_8_5_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10841 downto 10840)));
	track_8_5_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10843 downto 10842)));
	track_8_5_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10845 downto 10844)));
	track_8_5_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10847 downto 10846)));
	track_8_5_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10849 downto 10848)));
	track_8_5_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10851 downto 10850)));
	track_8_5_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10853 downto 10852)));
	track_8_5_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10855 downto 10854)));
	track_8_5_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10857 downto 10856)));
	track_8_5_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10859 downto 10858)));
	track_8_5_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10861 downto 10860)));
	track_8_5_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10863 downto 10862)));
	track_8_5_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10865 downto 10864)));
	track_8_5_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10867 downto 10866)));
	track_8_5_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10869 downto 10868)));
	track_8_5_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10871 downto 10870)));
	track_8_5_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10873 downto 10872)));
	track_8_5_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10875 downto 10874)));
	track_8_5_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10877 downto 10876)));
	track_8_5_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10879 downto 10878)));
	track_8_5_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10881 downto 10880)));
	track_8_5_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10883 downto 10882)));
	track_8_5_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10885 downto 10884)));
	track_8_5_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10887 downto 10886)));
	track_8_5_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10889 downto 10888)));
	track_8_5_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10891 downto 10890)));
	track_8_5_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10893 downto 10892)));
	track_8_5_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10895 downto 10894)));
	track_8_6_chanX_n0_driver_mux_selector  <= to_integer(unsigned(config(10897 downto 10896)));
	track_8_6_chanX_n1_driver_mux_selector  <= to_integer(unsigned(config(10899 downto 10898)));
	track_8_6_chanX_n10_driver_mux_selector <= to_integer(unsigned(config(10901 downto 10900)));
	track_8_6_chanX_n11_driver_mux_selector <= to_integer(unsigned(config(10902 downto 10902)));
	track_8_6_chanX_n12_driver_mux_selector <= to_integer(unsigned(config(10904 downto 10903)));
	track_8_6_chanX_n13_driver_mux_selector <= to_integer(unsigned(config(10905 downto 10905)));
	track_8_6_chanX_n14_driver_mux_selector <= to_integer(unsigned(config(10907 downto 10906)));
	track_8_6_chanX_n15_driver_mux_selector <= to_integer(unsigned(config(10908 downto 10908)));
	track_8_6_chanX_n2_driver_mux_selector  <= to_integer(unsigned(config(10910 downto 10909)));
	track_8_6_chanX_n3_driver_mux_selector  <= to_integer(unsigned(config(10912 downto 10911)));
	track_8_6_chanX_n4_driver_mux_selector  <= to_integer(unsigned(config(10914 downto 10913)));
	track_8_6_chanX_n5_driver_mux_selector  <= to_integer(unsigned(config(10916 downto 10915)));
	track_8_6_chanX_n6_driver_mux_selector  <= to_integer(unsigned(config(10918 downto 10917)));
	track_8_6_chanX_n7_driver_mux_selector  <= to_integer(unsigned(config(10920 downto 10919)));
	track_8_6_chanX_n8_driver_mux_selector  <= to_integer(unsigned(config(10922 downto 10921)));
	track_8_6_chanX_n9_driver_mux_selector  <= to_integer(unsigned(config(10923 downto 10923)));
	track_8_6_chanY_n0_driver_mux_selector  <= to_integer(unsigned(config(10925 downto 10924)));
	track_8_6_chanY_n1_driver_mux_selector  <= to_integer(unsigned(config(10927 downto 10926)));
	track_8_6_chanY_n10_driver_mux_selector <= to_integer(unsigned(config(10929 downto 10928)));
	track_8_6_chanY_n11_driver_mux_selector <= to_integer(unsigned(config(10930 downto 10930)));
	track_8_6_chanY_n12_driver_mux_selector <= to_integer(unsigned(config(10932 downto 10931)));
	track_8_6_chanY_n13_driver_mux_selector <= to_integer(unsigned(config(10933 downto 10933)));
	track_8_6_chanY_n14_driver_mux_selector <= to_integer(unsigned(config(10935 downto 10934)));
	track_8_6_chanY_n15_driver_mux_selector <= to_integer(unsigned(config(10936 downto 10936)));
	track_8_6_chanY_n2_driver_mux_selector  <= to_integer(unsigned(config(10938 downto 10937)));
	track_8_6_chanY_n3_driver_mux_selector  <= to_integer(unsigned(config(10940 downto 10939)));
	track_8_6_chanY_n4_driver_mux_selector  <= to_integer(unsigned(config(10942 downto 10941)));
	track_8_6_chanY_n5_driver_mux_selector  <= to_integer(unsigned(config(10944 downto 10943)));
	track_8_6_chanY_n6_driver_mux_selector  <= to_integer(unsigned(config(10946 downto 10945)));
	track_8_6_chanY_n7_driver_mux_selector  <= to_integer(unsigned(config(10948 downto 10947)));
	track_8_6_chanY_n8_driver_mux_selector  <= to_integer(unsigned(config(10950 downto 10949)));
	track_8_6_chanY_n9_driver_mux_selector  <= to_integer(unsigned(config(10951 downto 10951)));

	-- Tracks --
	-- All tracks are driven by a multiplexeur whose output is registered in a VTPR --
	process(clk)
	begin
		if rising_edge(clk) then
			track_0_1_chanY_n0  <= track_0_1_chanY_n0_driver_mux_fanins(track_0_1_chanY_n0_driver_mux_selector);
			track_0_1_chanY_n1  <= track_0_1_chanY_n1_driver_mux_fanins(track_0_1_chanY_n1_driver_mux_selector);
			track_0_1_chanY_n10 <= track_0_1_chanY_n10_driver_mux_fanins(track_0_1_chanY_n10_driver_mux_selector);
			track_0_1_chanY_n11 <= track_0_1_chanY_n11_driver_mux_fanins(track_0_1_chanY_n11_driver_mux_selector);
			track_0_1_chanY_n12 <= track_0_1_chanY_n12_driver_mux_fanins(track_0_1_chanY_n12_driver_mux_selector);
			track_0_1_chanY_n13 <= track_0_1_chanY_n13_driver_mux_fanins(track_0_1_chanY_n13_driver_mux_selector);
			track_0_1_chanY_n14 <= track_0_1_chanY_n14_driver_mux_fanins(track_0_1_chanY_n14_driver_mux_selector);
			track_0_1_chanY_n15 <= track_0_1_chanY_n15_driver_mux_fanins(track_0_1_chanY_n15_driver_mux_selector);
			track_0_1_chanY_n2  <= track_0_1_chanY_n2_driver_mux_fanins(track_0_1_chanY_n2_driver_mux_selector);
			track_0_1_chanY_n3  <= track_0_1_chanY_n3_driver_mux_fanins(track_0_1_chanY_n3_driver_mux_selector);
			track_0_1_chanY_n4  <= track_0_1_chanY_n4_driver_mux_fanins(track_0_1_chanY_n4_driver_mux_selector);
			track_0_1_chanY_n5  <= track_0_1_chanY_n5_driver_mux_fanins(track_0_1_chanY_n5_driver_mux_selector);
			track_0_1_chanY_n6  <= track_0_1_chanY_n6_driver_mux_fanins(track_0_1_chanY_n6_driver_mux_selector);
			track_0_1_chanY_n7  <= track_0_1_chanY_n7_driver_mux_fanins(track_0_1_chanY_n7_driver_mux_selector);
			track_0_1_chanY_n8  <= track_0_1_chanY_n8_driver_mux_fanins(track_0_1_chanY_n8_driver_mux_selector);
			track_0_1_chanY_n9  <= track_0_1_chanY_n9_driver_mux_fanins(track_0_1_chanY_n9_driver_mux_selector);
			track_0_2_chanY_n0  <= track_0_2_chanY_n0_driver_mux_fanins(track_0_2_chanY_n0_driver_mux_selector);
			track_0_2_chanY_n1  <= track_0_2_chanY_n1_driver_mux_fanins(track_0_2_chanY_n1_driver_mux_selector);
			track_0_2_chanY_n10 <= track_0_2_chanY_n10_driver_mux_fanins(track_0_2_chanY_n10_driver_mux_selector);
			track_0_2_chanY_n11 <= track_0_2_chanY_n11_driver_mux_fanins(track_0_2_chanY_n11_driver_mux_selector);
			track_0_2_chanY_n12 <= track_0_2_chanY_n12_driver_mux_fanins(track_0_2_chanY_n12_driver_mux_selector);
			track_0_2_chanY_n13 <= track_0_2_chanY_n13_driver_mux_fanins(track_0_2_chanY_n13_driver_mux_selector);
			track_0_2_chanY_n14 <= track_0_2_chanY_n14_driver_mux_fanins(track_0_2_chanY_n14_driver_mux_selector);
			track_0_2_chanY_n15 <= track_0_2_chanY_n15_driver_mux_fanins(track_0_2_chanY_n15_driver_mux_selector);
			track_0_2_chanY_n2  <= track_0_2_chanY_n2_driver_mux_fanins(track_0_2_chanY_n2_driver_mux_selector);
			track_0_2_chanY_n3  <= track_0_2_chanY_n3_driver_mux_fanins(track_0_2_chanY_n3_driver_mux_selector);
			track_0_2_chanY_n4  <= track_0_2_chanY_n4_driver_mux_fanins(track_0_2_chanY_n4_driver_mux_selector);
			track_0_2_chanY_n5  <= track_0_2_chanY_n5_driver_mux_fanins(track_0_2_chanY_n5_driver_mux_selector);
			track_0_2_chanY_n6  <= track_0_2_chanY_n6_driver_mux_fanins(track_0_2_chanY_n6_driver_mux_selector);
			track_0_2_chanY_n7  <= track_0_2_chanY_n7_driver_mux_fanins(track_0_2_chanY_n7_driver_mux_selector);
			track_0_2_chanY_n8  <= track_0_2_chanY_n8_driver_mux_fanins(track_0_2_chanY_n8_driver_mux_selector);
			track_0_2_chanY_n9  <= track_0_2_chanY_n9_driver_mux_fanins(track_0_2_chanY_n9_driver_mux_selector);
			track_0_3_chanY_n0  <= track_0_3_chanY_n0_driver_mux_fanins(track_0_3_chanY_n0_driver_mux_selector);
			track_0_3_chanY_n1  <= track_0_3_chanY_n1_driver_mux_fanins(track_0_3_chanY_n1_driver_mux_selector);
			track_0_3_chanY_n10 <= track_0_3_chanY_n10_driver_mux_fanins(track_0_3_chanY_n10_driver_mux_selector);
			track_0_3_chanY_n11 <= track_0_3_chanY_n11_driver_mux_fanins(track_0_3_chanY_n11_driver_mux_selector);
			track_0_3_chanY_n12 <= track_0_3_chanY_n12_driver_mux_fanins(track_0_3_chanY_n12_driver_mux_selector);
			track_0_3_chanY_n13 <= track_0_3_chanY_n13_driver_mux_fanins(track_0_3_chanY_n13_driver_mux_selector);
			track_0_3_chanY_n14 <= track_0_3_chanY_n14_driver_mux_fanins(track_0_3_chanY_n14_driver_mux_selector);
			track_0_3_chanY_n15 <= track_0_3_chanY_n15_driver_mux_fanins(track_0_3_chanY_n15_driver_mux_selector);
			track_0_3_chanY_n2  <= track_0_3_chanY_n2_driver_mux_fanins(track_0_3_chanY_n2_driver_mux_selector);
			track_0_3_chanY_n3  <= track_0_3_chanY_n3_driver_mux_fanins(track_0_3_chanY_n3_driver_mux_selector);
			track_0_3_chanY_n4  <= track_0_3_chanY_n4_driver_mux_fanins(track_0_3_chanY_n4_driver_mux_selector);
			track_0_3_chanY_n5  <= track_0_3_chanY_n5_driver_mux_fanins(track_0_3_chanY_n5_driver_mux_selector);
			track_0_3_chanY_n6  <= track_0_3_chanY_n6_driver_mux_fanins(track_0_3_chanY_n6_driver_mux_selector);
			track_0_3_chanY_n7  <= track_0_3_chanY_n7_driver_mux_fanins(track_0_3_chanY_n7_driver_mux_selector);
			track_0_3_chanY_n8  <= track_0_3_chanY_n8_driver_mux_fanins(track_0_3_chanY_n8_driver_mux_selector);
			track_0_3_chanY_n9  <= track_0_3_chanY_n9_driver_mux_fanins(track_0_3_chanY_n9_driver_mux_selector);
			track_0_4_chanY_n0  <= track_0_4_chanY_n0_driver_mux_fanins(track_0_4_chanY_n0_driver_mux_selector);
			track_0_4_chanY_n1  <= track_0_4_chanY_n1_driver_mux_fanins(track_0_4_chanY_n1_driver_mux_selector);
			track_0_4_chanY_n10 <= track_0_4_chanY_n10_driver_mux_fanins(track_0_4_chanY_n10_driver_mux_selector);
			track_0_4_chanY_n11 <= track_0_4_chanY_n11_driver_mux_fanins(track_0_4_chanY_n11_driver_mux_selector);
			track_0_4_chanY_n12 <= track_0_4_chanY_n12_driver_mux_fanins(track_0_4_chanY_n12_driver_mux_selector);
			track_0_4_chanY_n13 <= track_0_4_chanY_n13_driver_mux_fanins(track_0_4_chanY_n13_driver_mux_selector);
			track_0_4_chanY_n14 <= track_0_4_chanY_n14_driver_mux_fanins(track_0_4_chanY_n14_driver_mux_selector);
			track_0_4_chanY_n15 <= track_0_4_chanY_n15_driver_mux_fanins(track_0_4_chanY_n15_driver_mux_selector);
			track_0_4_chanY_n2  <= track_0_4_chanY_n2_driver_mux_fanins(track_0_4_chanY_n2_driver_mux_selector);
			track_0_4_chanY_n3  <= track_0_4_chanY_n3_driver_mux_fanins(track_0_4_chanY_n3_driver_mux_selector);
			track_0_4_chanY_n4  <= track_0_4_chanY_n4_driver_mux_fanins(track_0_4_chanY_n4_driver_mux_selector);
			track_0_4_chanY_n5  <= track_0_4_chanY_n5_driver_mux_fanins(track_0_4_chanY_n5_driver_mux_selector);
			track_0_4_chanY_n6  <= track_0_4_chanY_n6_driver_mux_fanins(track_0_4_chanY_n6_driver_mux_selector);
			track_0_4_chanY_n7  <= track_0_4_chanY_n7_driver_mux_fanins(track_0_4_chanY_n7_driver_mux_selector);
			track_0_4_chanY_n8  <= track_0_4_chanY_n8_driver_mux_fanins(track_0_4_chanY_n8_driver_mux_selector);
			track_0_4_chanY_n9  <= track_0_4_chanY_n9_driver_mux_fanins(track_0_4_chanY_n9_driver_mux_selector);
			track_0_5_chanY_n0  <= track_0_5_chanY_n0_driver_mux_fanins(track_0_5_chanY_n0_driver_mux_selector);
			track_0_5_chanY_n1  <= track_0_5_chanY_n1_driver_mux_fanins(track_0_5_chanY_n1_driver_mux_selector);
			track_0_5_chanY_n10 <= track_0_5_chanY_n10_driver_mux_fanins(track_0_5_chanY_n10_driver_mux_selector);
			track_0_5_chanY_n11 <= track_0_5_chanY_n11_driver_mux_fanins(track_0_5_chanY_n11_driver_mux_selector);
			track_0_5_chanY_n12 <= track_0_5_chanY_n12_driver_mux_fanins(track_0_5_chanY_n12_driver_mux_selector);
			track_0_5_chanY_n13 <= track_0_5_chanY_n13_driver_mux_fanins(track_0_5_chanY_n13_driver_mux_selector);
			track_0_5_chanY_n14 <= track_0_5_chanY_n14_driver_mux_fanins(track_0_5_chanY_n14_driver_mux_selector);
			track_0_5_chanY_n15 <= track_0_5_chanY_n15_driver_mux_fanins(track_0_5_chanY_n15_driver_mux_selector);
			track_0_5_chanY_n2  <= track_0_5_chanY_n2_driver_mux_fanins(track_0_5_chanY_n2_driver_mux_selector);
			track_0_5_chanY_n3  <= track_0_5_chanY_n3_driver_mux_fanins(track_0_5_chanY_n3_driver_mux_selector);
			track_0_5_chanY_n4  <= track_0_5_chanY_n4_driver_mux_fanins(track_0_5_chanY_n4_driver_mux_selector);
			track_0_5_chanY_n5  <= track_0_5_chanY_n5_driver_mux_fanins(track_0_5_chanY_n5_driver_mux_selector);
			track_0_5_chanY_n6  <= track_0_5_chanY_n6_driver_mux_fanins(track_0_5_chanY_n6_driver_mux_selector);
			track_0_5_chanY_n7  <= track_0_5_chanY_n7_driver_mux_fanins(track_0_5_chanY_n7_driver_mux_selector);
			track_0_5_chanY_n8  <= track_0_5_chanY_n8_driver_mux_fanins(track_0_5_chanY_n8_driver_mux_selector);
			track_0_5_chanY_n9  <= track_0_5_chanY_n9_driver_mux_fanins(track_0_5_chanY_n9_driver_mux_selector);
			track_0_6_chanY_n0  <= track_0_6_chanY_n0_driver_mux_fanins(track_0_6_chanY_n0_driver_mux_selector);
			track_0_6_chanY_n1  <= track_0_6_chanY_n1_driver_mux_fanins(track_0_6_chanY_n1_driver_mux_selector);
			track_0_6_chanY_n10 <= track_0_6_chanY_n10_driver_mux_fanins(track_0_6_chanY_n10_driver_mux_selector);
			track_0_6_chanY_n11 <= track_0_6_chanY_n11_driver_mux_fanins(track_0_6_chanY_n11_driver_mux_selector);
			track_0_6_chanY_n12 <= track_0_6_chanY_n12_driver_mux_fanins(track_0_6_chanY_n12_driver_mux_selector);
			track_0_6_chanY_n13 <= track_0_6_chanY_n13_driver_mux_fanins(track_0_6_chanY_n13_driver_mux_selector);
			track_0_6_chanY_n14 <= track_0_6_chanY_n14_driver_mux_fanins(track_0_6_chanY_n14_driver_mux_selector);
			track_0_6_chanY_n15 <= track_0_6_chanY_n15_driver_mux_fanins(track_0_6_chanY_n15_driver_mux_selector);
			track_0_6_chanY_n2  <= track_0_6_chanY_n2_driver_mux_fanins(track_0_6_chanY_n2_driver_mux_selector);
			track_0_6_chanY_n3  <= track_0_6_chanY_n3_driver_mux_fanins(track_0_6_chanY_n3_driver_mux_selector);
			track_0_6_chanY_n4  <= track_0_6_chanY_n4_driver_mux_fanins(track_0_6_chanY_n4_driver_mux_selector);
			track_0_6_chanY_n5  <= track_0_6_chanY_n5_driver_mux_fanins(track_0_6_chanY_n5_driver_mux_selector);
			track_0_6_chanY_n6  <= track_0_6_chanY_n6_driver_mux_fanins(track_0_6_chanY_n6_driver_mux_selector);
			track_0_6_chanY_n7  <= track_0_6_chanY_n7_driver_mux_fanins(track_0_6_chanY_n7_driver_mux_selector);
			track_0_6_chanY_n8  <= track_0_6_chanY_n8_driver_mux_fanins(track_0_6_chanY_n8_driver_mux_selector);
			track_0_6_chanY_n9  <= track_0_6_chanY_n9_driver_mux_fanins(track_0_6_chanY_n9_driver_mux_selector);
			track_1_0_chanX_n0  <= track_1_0_chanX_n0_driver_mux_fanins(track_1_0_chanX_n0_driver_mux_selector);
			track_1_0_chanX_n1  <= track_1_0_chanX_n1_driver_mux_fanins(track_1_0_chanX_n1_driver_mux_selector);
			track_1_0_chanX_n10 <= track_1_0_chanX_n10_driver_mux_fanins(track_1_0_chanX_n10_driver_mux_selector);
			track_1_0_chanX_n11 <= track_1_0_chanX_n11_driver_mux_fanins(track_1_0_chanX_n11_driver_mux_selector);
			track_1_0_chanX_n12 <= track_1_0_chanX_n12_driver_mux_fanins(track_1_0_chanX_n12_driver_mux_selector);
			track_1_0_chanX_n13 <= track_1_0_chanX_n13_driver_mux_fanins(track_1_0_chanX_n13_driver_mux_selector);
			track_1_0_chanX_n14 <= track_1_0_chanX_n14_driver_mux_fanins(track_1_0_chanX_n14_driver_mux_selector);
			track_1_0_chanX_n15 <= track_1_0_chanX_n15_driver_mux_fanins(track_1_0_chanX_n15_driver_mux_selector);
			track_1_0_chanX_n2  <= track_1_0_chanX_n2_driver_mux_fanins(track_1_0_chanX_n2_driver_mux_selector);
			track_1_0_chanX_n3  <= track_1_0_chanX_n3_driver_mux_fanins(track_1_0_chanX_n3_driver_mux_selector);
			track_1_0_chanX_n4  <= track_1_0_chanX_n4_driver_mux_fanins(track_1_0_chanX_n4_driver_mux_selector);
			track_1_0_chanX_n5  <= track_1_0_chanX_n5_driver_mux_fanins(track_1_0_chanX_n5_driver_mux_selector);
			track_1_0_chanX_n6  <= track_1_0_chanX_n6_driver_mux_fanins(track_1_0_chanX_n6_driver_mux_selector);
			track_1_0_chanX_n7  <= track_1_0_chanX_n7_driver_mux_fanins(track_1_0_chanX_n7_driver_mux_selector);
			track_1_0_chanX_n8  <= track_1_0_chanX_n8_driver_mux_fanins(track_1_0_chanX_n8_driver_mux_selector);
			track_1_0_chanX_n9  <= track_1_0_chanX_n9_driver_mux_fanins(track_1_0_chanX_n9_driver_mux_selector);
			track_1_1_chanX_n0  <= track_1_1_chanX_n0_driver_mux_fanins(track_1_1_chanX_n0_driver_mux_selector);
			track_1_1_chanX_n1  <= track_1_1_chanX_n1_driver_mux_fanins(track_1_1_chanX_n1_driver_mux_selector);
			track_1_1_chanX_n10 <= track_1_1_chanX_n10_driver_mux_fanins(track_1_1_chanX_n10_driver_mux_selector);
			track_1_1_chanX_n11 <= track_1_1_chanX_n11_driver_mux_fanins(track_1_1_chanX_n11_driver_mux_selector);
			track_1_1_chanX_n12 <= track_1_1_chanX_n12_driver_mux_fanins(track_1_1_chanX_n12_driver_mux_selector);
			track_1_1_chanX_n13 <= track_1_1_chanX_n13_driver_mux_fanins(track_1_1_chanX_n13_driver_mux_selector);
			track_1_1_chanX_n14 <= track_1_1_chanX_n14_driver_mux_fanins(track_1_1_chanX_n14_driver_mux_selector);
			track_1_1_chanX_n15 <= track_1_1_chanX_n15_driver_mux_fanins(track_1_1_chanX_n15_driver_mux_selector);
			track_1_1_chanX_n2  <= track_1_1_chanX_n2_driver_mux_fanins(track_1_1_chanX_n2_driver_mux_selector);
			track_1_1_chanX_n3  <= track_1_1_chanX_n3_driver_mux_fanins(track_1_1_chanX_n3_driver_mux_selector);
			track_1_1_chanX_n4  <= track_1_1_chanX_n4_driver_mux_fanins(track_1_1_chanX_n4_driver_mux_selector);
			track_1_1_chanX_n5  <= track_1_1_chanX_n5_driver_mux_fanins(track_1_1_chanX_n5_driver_mux_selector);
			track_1_1_chanX_n6  <= track_1_1_chanX_n6_driver_mux_fanins(track_1_1_chanX_n6_driver_mux_selector);
			track_1_1_chanX_n7  <= track_1_1_chanX_n7_driver_mux_fanins(track_1_1_chanX_n7_driver_mux_selector);
			track_1_1_chanX_n8  <= track_1_1_chanX_n8_driver_mux_fanins(track_1_1_chanX_n8_driver_mux_selector);
			track_1_1_chanX_n9  <= track_1_1_chanX_n9_driver_mux_fanins(track_1_1_chanX_n9_driver_mux_selector);
			track_1_1_chanY_n0  <= track_1_1_chanY_n0_driver_mux_fanins(track_1_1_chanY_n0_driver_mux_selector);
			track_1_1_chanY_n1  <= track_1_1_chanY_n1_driver_mux_fanins(track_1_1_chanY_n1_driver_mux_selector);
			track_1_1_chanY_n10 <= track_1_1_chanY_n10_driver_mux_fanins(track_1_1_chanY_n10_driver_mux_selector);
			track_1_1_chanY_n11 <= track_1_1_chanY_n11_driver_mux_fanins(track_1_1_chanY_n11_driver_mux_selector);
			track_1_1_chanY_n12 <= track_1_1_chanY_n12_driver_mux_fanins(track_1_1_chanY_n12_driver_mux_selector);
			track_1_1_chanY_n13 <= track_1_1_chanY_n13_driver_mux_fanins(track_1_1_chanY_n13_driver_mux_selector);
			track_1_1_chanY_n14 <= track_1_1_chanY_n14_driver_mux_fanins(track_1_1_chanY_n14_driver_mux_selector);
			track_1_1_chanY_n15 <= track_1_1_chanY_n15_driver_mux_fanins(track_1_1_chanY_n15_driver_mux_selector);
			track_1_1_chanY_n2  <= track_1_1_chanY_n2_driver_mux_fanins(track_1_1_chanY_n2_driver_mux_selector);
			track_1_1_chanY_n3  <= track_1_1_chanY_n3_driver_mux_fanins(track_1_1_chanY_n3_driver_mux_selector);
			track_1_1_chanY_n4  <= track_1_1_chanY_n4_driver_mux_fanins(track_1_1_chanY_n4_driver_mux_selector);
			track_1_1_chanY_n5  <= track_1_1_chanY_n5_driver_mux_fanins(track_1_1_chanY_n5_driver_mux_selector);
			track_1_1_chanY_n6  <= track_1_1_chanY_n6_driver_mux_fanins(track_1_1_chanY_n6_driver_mux_selector);
			track_1_1_chanY_n7  <= track_1_1_chanY_n7_driver_mux_fanins(track_1_1_chanY_n7_driver_mux_selector);
			track_1_1_chanY_n8  <= track_1_1_chanY_n8_driver_mux_fanins(track_1_1_chanY_n8_driver_mux_selector);
			track_1_1_chanY_n9  <= track_1_1_chanY_n9_driver_mux_fanins(track_1_1_chanY_n9_driver_mux_selector);
			track_1_2_chanX_n0  <= track_1_2_chanX_n0_driver_mux_fanins(track_1_2_chanX_n0_driver_mux_selector);
			track_1_2_chanX_n1  <= track_1_2_chanX_n1_driver_mux_fanins(track_1_2_chanX_n1_driver_mux_selector);
			track_1_2_chanX_n10 <= track_1_2_chanX_n10_driver_mux_fanins(track_1_2_chanX_n10_driver_mux_selector);
			track_1_2_chanX_n11 <= track_1_2_chanX_n11_driver_mux_fanins(track_1_2_chanX_n11_driver_mux_selector);
			track_1_2_chanX_n12 <= track_1_2_chanX_n12_driver_mux_fanins(track_1_2_chanX_n12_driver_mux_selector);
			track_1_2_chanX_n13 <= track_1_2_chanX_n13_driver_mux_fanins(track_1_2_chanX_n13_driver_mux_selector);
			track_1_2_chanX_n14 <= track_1_2_chanX_n14_driver_mux_fanins(track_1_2_chanX_n14_driver_mux_selector);
			track_1_2_chanX_n15 <= track_1_2_chanX_n15_driver_mux_fanins(track_1_2_chanX_n15_driver_mux_selector);
			track_1_2_chanX_n2  <= track_1_2_chanX_n2_driver_mux_fanins(track_1_2_chanX_n2_driver_mux_selector);
			track_1_2_chanX_n3  <= track_1_2_chanX_n3_driver_mux_fanins(track_1_2_chanX_n3_driver_mux_selector);
			track_1_2_chanX_n4  <= track_1_2_chanX_n4_driver_mux_fanins(track_1_2_chanX_n4_driver_mux_selector);
			track_1_2_chanX_n5  <= track_1_2_chanX_n5_driver_mux_fanins(track_1_2_chanX_n5_driver_mux_selector);
			track_1_2_chanX_n6  <= track_1_2_chanX_n6_driver_mux_fanins(track_1_2_chanX_n6_driver_mux_selector);
			track_1_2_chanX_n7  <= track_1_2_chanX_n7_driver_mux_fanins(track_1_2_chanX_n7_driver_mux_selector);
			track_1_2_chanX_n8  <= track_1_2_chanX_n8_driver_mux_fanins(track_1_2_chanX_n8_driver_mux_selector);
			track_1_2_chanX_n9  <= track_1_2_chanX_n9_driver_mux_fanins(track_1_2_chanX_n9_driver_mux_selector);
			track_1_2_chanY_n0  <= track_1_2_chanY_n0_driver_mux_fanins(track_1_2_chanY_n0_driver_mux_selector);
			track_1_2_chanY_n1  <= track_1_2_chanY_n1_driver_mux_fanins(track_1_2_chanY_n1_driver_mux_selector);
			track_1_2_chanY_n10 <= track_1_2_chanY_n10_driver_mux_fanins(track_1_2_chanY_n10_driver_mux_selector);
			track_1_2_chanY_n11 <= track_1_2_chanY_n11_driver_mux_fanins(track_1_2_chanY_n11_driver_mux_selector);
			track_1_2_chanY_n12 <= track_1_2_chanY_n12_driver_mux_fanins(track_1_2_chanY_n12_driver_mux_selector);
			track_1_2_chanY_n13 <= track_1_2_chanY_n13_driver_mux_fanins(track_1_2_chanY_n13_driver_mux_selector);
			track_1_2_chanY_n14 <= track_1_2_chanY_n14_driver_mux_fanins(track_1_2_chanY_n14_driver_mux_selector);
			track_1_2_chanY_n15 <= track_1_2_chanY_n15_driver_mux_fanins(track_1_2_chanY_n15_driver_mux_selector);
			track_1_2_chanY_n2  <= track_1_2_chanY_n2_driver_mux_fanins(track_1_2_chanY_n2_driver_mux_selector);
			track_1_2_chanY_n3  <= track_1_2_chanY_n3_driver_mux_fanins(track_1_2_chanY_n3_driver_mux_selector);
			track_1_2_chanY_n4  <= track_1_2_chanY_n4_driver_mux_fanins(track_1_2_chanY_n4_driver_mux_selector);
			track_1_2_chanY_n5  <= track_1_2_chanY_n5_driver_mux_fanins(track_1_2_chanY_n5_driver_mux_selector);
			track_1_2_chanY_n6  <= track_1_2_chanY_n6_driver_mux_fanins(track_1_2_chanY_n6_driver_mux_selector);
			track_1_2_chanY_n7  <= track_1_2_chanY_n7_driver_mux_fanins(track_1_2_chanY_n7_driver_mux_selector);
			track_1_2_chanY_n8  <= track_1_2_chanY_n8_driver_mux_fanins(track_1_2_chanY_n8_driver_mux_selector);
			track_1_2_chanY_n9  <= track_1_2_chanY_n9_driver_mux_fanins(track_1_2_chanY_n9_driver_mux_selector);
			track_1_3_chanX_n0  <= track_1_3_chanX_n0_driver_mux_fanins(track_1_3_chanX_n0_driver_mux_selector);
			track_1_3_chanX_n1  <= track_1_3_chanX_n1_driver_mux_fanins(track_1_3_chanX_n1_driver_mux_selector);
			track_1_3_chanX_n10 <= track_1_3_chanX_n10_driver_mux_fanins(track_1_3_chanX_n10_driver_mux_selector);
			track_1_3_chanX_n11 <= track_1_3_chanX_n11_driver_mux_fanins(track_1_3_chanX_n11_driver_mux_selector);
			track_1_3_chanX_n12 <= track_1_3_chanX_n12_driver_mux_fanins(track_1_3_chanX_n12_driver_mux_selector);
			track_1_3_chanX_n13 <= track_1_3_chanX_n13_driver_mux_fanins(track_1_3_chanX_n13_driver_mux_selector);
			track_1_3_chanX_n14 <= track_1_3_chanX_n14_driver_mux_fanins(track_1_3_chanX_n14_driver_mux_selector);
			track_1_3_chanX_n15 <= track_1_3_chanX_n15_driver_mux_fanins(track_1_3_chanX_n15_driver_mux_selector);
			track_1_3_chanX_n2  <= track_1_3_chanX_n2_driver_mux_fanins(track_1_3_chanX_n2_driver_mux_selector);
			track_1_3_chanX_n3  <= track_1_3_chanX_n3_driver_mux_fanins(track_1_3_chanX_n3_driver_mux_selector);
			track_1_3_chanX_n4  <= track_1_3_chanX_n4_driver_mux_fanins(track_1_3_chanX_n4_driver_mux_selector);
			track_1_3_chanX_n5  <= track_1_3_chanX_n5_driver_mux_fanins(track_1_3_chanX_n5_driver_mux_selector);
			track_1_3_chanX_n6  <= track_1_3_chanX_n6_driver_mux_fanins(track_1_3_chanX_n6_driver_mux_selector);
			track_1_3_chanX_n7  <= track_1_3_chanX_n7_driver_mux_fanins(track_1_3_chanX_n7_driver_mux_selector);
			track_1_3_chanX_n8  <= track_1_3_chanX_n8_driver_mux_fanins(track_1_3_chanX_n8_driver_mux_selector);
			track_1_3_chanX_n9  <= track_1_3_chanX_n9_driver_mux_fanins(track_1_3_chanX_n9_driver_mux_selector);
			track_1_3_chanY_n0  <= track_1_3_chanY_n0_driver_mux_fanins(track_1_3_chanY_n0_driver_mux_selector);
			track_1_3_chanY_n1  <= track_1_3_chanY_n1_driver_mux_fanins(track_1_3_chanY_n1_driver_mux_selector);
			track_1_3_chanY_n10 <= track_1_3_chanY_n10_driver_mux_fanins(track_1_3_chanY_n10_driver_mux_selector);
			track_1_3_chanY_n11 <= track_1_3_chanY_n11_driver_mux_fanins(track_1_3_chanY_n11_driver_mux_selector);
			track_1_3_chanY_n12 <= track_1_3_chanY_n12_driver_mux_fanins(track_1_3_chanY_n12_driver_mux_selector);
			track_1_3_chanY_n13 <= track_1_3_chanY_n13_driver_mux_fanins(track_1_3_chanY_n13_driver_mux_selector);
			track_1_3_chanY_n14 <= track_1_3_chanY_n14_driver_mux_fanins(track_1_3_chanY_n14_driver_mux_selector);
			track_1_3_chanY_n15 <= track_1_3_chanY_n15_driver_mux_fanins(track_1_3_chanY_n15_driver_mux_selector);
			track_1_3_chanY_n2  <= track_1_3_chanY_n2_driver_mux_fanins(track_1_3_chanY_n2_driver_mux_selector);
			track_1_3_chanY_n3  <= track_1_3_chanY_n3_driver_mux_fanins(track_1_3_chanY_n3_driver_mux_selector);
			track_1_3_chanY_n4  <= track_1_3_chanY_n4_driver_mux_fanins(track_1_3_chanY_n4_driver_mux_selector);
			track_1_3_chanY_n5  <= track_1_3_chanY_n5_driver_mux_fanins(track_1_3_chanY_n5_driver_mux_selector);
			track_1_3_chanY_n6  <= track_1_3_chanY_n6_driver_mux_fanins(track_1_3_chanY_n6_driver_mux_selector);
			track_1_3_chanY_n7  <= track_1_3_chanY_n7_driver_mux_fanins(track_1_3_chanY_n7_driver_mux_selector);
			track_1_3_chanY_n8  <= track_1_3_chanY_n8_driver_mux_fanins(track_1_3_chanY_n8_driver_mux_selector);
			track_1_3_chanY_n9  <= track_1_3_chanY_n9_driver_mux_fanins(track_1_3_chanY_n9_driver_mux_selector);
			track_1_4_chanX_n0  <= track_1_4_chanX_n0_driver_mux_fanins(track_1_4_chanX_n0_driver_mux_selector);
			track_1_4_chanX_n1  <= track_1_4_chanX_n1_driver_mux_fanins(track_1_4_chanX_n1_driver_mux_selector);
			track_1_4_chanX_n10 <= track_1_4_chanX_n10_driver_mux_fanins(track_1_4_chanX_n10_driver_mux_selector);
			track_1_4_chanX_n11 <= track_1_4_chanX_n11_driver_mux_fanins(track_1_4_chanX_n11_driver_mux_selector);
			track_1_4_chanX_n12 <= track_1_4_chanX_n12_driver_mux_fanins(track_1_4_chanX_n12_driver_mux_selector);
			track_1_4_chanX_n13 <= track_1_4_chanX_n13_driver_mux_fanins(track_1_4_chanX_n13_driver_mux_selector);
			track_1_4_chanX_n14 <= track_1_4_chanX_n14_driver_mux_fanins(track_1_4_chanX_n14_driver_mux_selector);
			track_1_4_chanX_n15 <= track_1_4_chanX_n15_driver_mux_fanins(track_1_4_chanX_n15_driver_mux_selector);
			track_1_4_chanX_n2  <= track_1_4_chanX_n2_driver_mux_fanins(track_1_4_chanX_n2_driver_mux_selector);
			track_1_4_chanX_n3  <= track_1_4_chanX_n3_driver_mux_fanins(track_1_4_chanX_n3_driver_mux_selector);
			track_1_4_chanX_n4  <= track_1_4_chanX_n4_driver_mux_fanins(track_1_4_chanX_n4_driver_mux_selector);
			track_1_4_chanX_n5  <= track_1_4_chanX_n5_driver_mux_fanins(track_1_4_chanX_n5_driver_mux_selector);
			track_1_4_chanX_n6  <= track_1_4_chanX_n6_driver_mux_fanins(track_1_4_chanX_n6_driver_mux_selector);
			track_1_4_chanX_n7  <= track_1_4_chanX_n7_driver_mux_fanins(track_1_4_chanX_n7_driver_mux_selector);
			track_1_4_chanX_n8  <= track_1_4_chanX_n8_driver_mux_fanins(track_1_4_chanX_n8_driver_mux_selector);
			track_1_4_chanX_n9  <= track_1_4_chanX_n9_driver_mux_fanins(track_1_4_chanX_n9_driver_mux_selector);
			track_1_4_chanY_n0  <= track_1_4_chanY_n0_driver_mux_fanins(track_1_4_chanY_n0_driver_mux_selector);
			track_1_4_chanY_n1  <= track_1_4_chanY_n1_driver_mux_fanins(track_1_4_chanY_n1_driver_mux_selector);
			track_1_4_chanY_n10 <= track_1_4_chanY_n10_driver_mux_fanins(track_1_4_chanY_n10_driver_mux_selector);
			track_1_4_chanY_n11 <= track_1_4_chanY_n11_driver_mux_fanins(track_1_4_chanY_n11_driver_mux_selector);
			track_1_4_chanY_n12 <= track_1_4_chanY_n12_driver_mux_fanins(track_1_4_chanY_n12_driver_mux_selector);
			track_1_4_chanY_n13 <= track_1_4_chanY_n13_driver_mux_fanins(track_1_4_chanY_n13_driver_mux_selector);
			track_1_4_chanY_n14 <= track_1_4_chanY_n14_driver_mux_fanins(track_1_4_chanY_n14_driver_mux_selector);
			track_1_4_chanY_n15 <= track_1_4_chanY_n15_driver_mux_fanins(track_1_4_chanY_n15_driver_mux_selector);
			track_1_4_chanY_n2  <= track_1_4_chanY_n2_driver_mux_fanins(track_1_4_chanY_n2_driver_mux_selector);
			track_1_4_chanY_n3  <= track_1_4_chanY_n3_driver_mux_fanins(track_1_4_chanY_n3_driver_mux_selector);
			track_1_4_chanY_n4  <= track_1_4_chanY_n4_driver_mux_fanins(track_1_4_chanY_n4_driver_mux_selector);
			track_1_4_chanY_n5  <= track_1_4_chanY_n5_driver_mux_fanins(track_1_4_chanY_n5_driver_mux_selector);
			track_1_4_chanY_n6  <= track_1_4_chanY_n6_driver_mux_fanins(track_1_4_chanY_n6_driver_mux_selector);
			track_1_4_chanY_n7  <= track_1_4_chanY_n7_driver_mux_fanins(track_1_4_chanY_n7_driver_mux_selector);
			track_1_4_chanY_n8  <= track_1_4_chanY_n8_driver_mux_fanins(track_1_4_chanY_n8_driver_mux_selector);
			track_1_4_chanY_n9  <= track_1_4_chanY_n9_driver_mux_fanins(track_1_4_chanY_n9_driver_mux_selector);
			track_1_5_chanX_n0  <= track_1_5_chanX_n0_driver_mux_fanins(track_1_5_chanX_n0_driver_mux_selector);
			track_1_5_chanX_n1  <= track_1_5_chanX_n1_driver_mux_fanins(track_1_5_chanX_n1_driver_mux_selector);
			track_1_5_chanX_n10 <= track_1_5_chanX_n10_driver_mux_fanins(track_1_5_chanX_n10_driver_mux_selector);
			track_1_5_chanX_n11 <= track_1_5_chanX_n11_driver_mux_fanins(track_1_5_chanX_n11_driver_mux_selector);
			track_1_5_chanX_n12 <= track_1_5_chanX_n12_driver_mux_fanins(track_1_5_chanX_n12_driver_mux_selector);
			track_1_5_chanX_n13 <= track_1_5_chanX_n13_driver_mux_fanins(track_1_5_chanX_n13_driver_mux_selector);
			track_1_5_chanX_n14 <= track_1_5_chanX_n14_driver_mux_fanins(track_1_5_chanX_n14_driver_mux_selector);
			track_1_5_chanX_n15 <= track_1_5_chanX_n15_driver_mux_fanins(track_1_5_chanX_n15_driver_mux_selector);
			track_1_5_chanX_n2  <= track_1_5_chanX_n2_driver_mux_fanins(track_1_5_chanX_n2_driver_mux_selector);
			track_1_5_chanX_n3  <= track_1_5_chanX_n3_driver_mux_fanins(track_1_5_chanX_n3_driver_mux_selector);
			track_1_5_chanX_n4  <= track_1_5_chanX_n4_driver_mux_fanins(track_1_5_chanX_n4_driver_mux_selector);
			track_1_5_chanX_n5  <= track_1_5_chanX_n5_driver_mux_fanins(track_1_5_chanX_n5_driver_mux_selector);
			track_1_5_chanX_n6  <= track_1_5_chanX_n6_driver_mux_fanins(track_1_5_chanX_n6_driver_mux_selector);
			track_1_5_chanX_n7  <= track_1_5_chanX_n7_driver_mux_fanins(track_1_5_chanX_n7_driver_mux_selector);
			track_1_5_chanX_n8  <= track_1_5_chanX_n8_driver_mux_fanins(track_1_5_chanX_n8_driver_mux_selector);
			track_1_5_chanX_n9  <= track_1_5_chanX_n9_driver_mux_fanins(track_1_5_chanX_n9_driver_mux_selector);
			track_1_5_chanY_n0  <= track_1_5_chanY_n0_driver_mux_fanins(track_1_5_chanY_n0_driver_mux_selector);
			track_1_5_chanY_n1  <= track_1_5_chanY_n1_driver_mux_fanins(track_1_5_chanY_n1_driver_mux_selector);
			track_1_5_chanY_n10 <= track_1_5_chanY_n10_driver_mux_fanins(track_1_5_chanY_n10_driver_mux_selector);
			track_1_5_chanY_n11 <= track_1_5_chanY_n11_driver_mux_fanins(track_1_5_chanY_n11_driver_mux_selector);
			track_1_5_chanY_n12 <= track_1_5_chanY_n12_driver_mux_fanins(track_1_5_chanY_n12_driver_mux_selector);
			track_1_5_chanY_n13 <= track_1_5_chanY_n13_driver_mux_fanins(track_1_5_chanY_n13_driver_mux_selector);
			track_1_5_chanY_n14 <= track_1_5_chanY_n14_driver_mux_fanins(track_1_5_chanY_n14_driver_mux_selector);
			track_1_5_chanY_n15 <= track_1_5_chanY_n15_driver_mux_fanins(track_1_5_chanY_n15_driver_mux_selector);
			track_1_5_chanY_n2  <= track_1_5_chanY_n2_driver_mux_fanins(track_1_5_chanY_n2_driver_mux_selector);
			track_1_5_chanY_n3  <= track_1_5_chanY_n3_driver_mux_fanins(track_1_5_chanY_n3_driver_mux_selector);
			track_1_5_chanY_n4  <= track_1_5_chanY_n4_driver_mux_fanins(track_1_5_chanY_n4_driver_mux_selector);
			track_1_5_chanY_n5  <= track_1_5_chanY_n5_driver_mux_fanins(track_1_5_chanY_n5_driver_mux_selector);
			track_1_5_chanY_n6  <= track_1_5_chanY_n6_driver_mux_fanins(track_1_5_chanY_n6_driver_mux_selector);
			track_1_5_chanY_n7  <= track_1_5_chanY_n7_driver_mux_fanins(track_1_5_chanY_n7_driver_mux_selector);
			track_1_5_chanY_n8  <= track_1_5_chanY_n8_driver_mux_fanins(track_1_5_chanY_n8_driver_mux_selector);
			track_1_5_chanY_n9  <= track_1_5_chanY_n9_driver_mux_fanins(track_1_5_chanY_n9_driver_mux_selector);
			track_1_6_chanX_n0  <= track_1_6_chanX_n0_driver_mux_fanins(track_1_6_chanX_n0_driver_mux_selector);
			track_1_6_chanX_n1  <= track_1_6_chanX_n1_driver_mux_fanins(track_1_6_chanX_n1_driver_mux_selector);
			track_1_6_chanX_n10 <= track_1_6_chanX_n10_driver_mux_fanins(track_1_6_chanX_n10_driver_mux_selector);
			track_1_6_chanX_n11 <= track_1_6_chanX_n11_driver_mux_fanins(track_1_6_chanX_n11_driver_mux_selector);
			track_1_6_chanX_n12 <= track_1_6_chanX_n12_driver_mux_fanins(track_1_6_chanX_n12_driver_mux_selector);
			track_1_6_chanX_n13 <= track_1_6_chanX_n13_driver_mux_fanins(track_1_6_chanX_n13_driver_mux_selector);
			track_1_6_chanX_n14 <= track_1_6_chanX_n14_driver_mux_fanins(track_1_6_chanX_n14_driver_mux_selector);
			track_1_6_chanX_n15 <= track_1_6_chanX_n15_driver_mux_fanins(track_1_6_chanX_n15_driver_mux_selector);
			track_1_6_chanX_n2  <= track_1_6_chanX_n2_driver_mux_fanins(track_1_6_chanX_n2_driver_mux_selector);
			track_1_6_chanX_n3  <= track_1_6_chanX_n3_driver_mux_fanins(track_1_6_chanX_n3_driver_mux_selector);
			track_1_6_chanX_n4  <= track_1_6_chanX_n4_driver_mux_fanins(track_1_6_chanX_n4_driver_mux_selector);
			track_1_6_chanX_n5  <= track_1_6_chanX_n5_driver_mux_fanins(track_1_6_chanX_n5_driver_mux_selector);
			track_1_6_chanX_n6  <= track_1_6_chanX_n6_driver_mux_fanins(track_1_6_chanX_n6_driver_mux_selector);
			track_1_6_chanX_n7  <= track_1_6_chanX_n7_driver_mux_fanins(track_1_6_chanX_n7_driver_mux_selector);
			track_1_6_chanX_n8  <= track_1_6_chanX_n8_driver_mux_fanins(track_1_6_chanX_n8_driver_mux_selector);
			track_1_6_chanX_n9  <= track_1_6_chanX_n9_driver_mux_fanins(track_1_6_chanX_n9_driver_mux_selector);
			track_1_6_chanY_n0  <= track_1_6_chanY_n0_driver_mux_fanins(track_1_6_chanY_n0_driver_mux_selector);
			track_1_6_chanY_n1  <= track_1_6_chanY_n1_driver_mux_fanins(track_1_6_chanY_n1_driver_mux_selector);
			track_1_6_chanY_n10 <= track_1_6_chanY_n10_driver_mux_fanins(track_1_6_chanY_n10_driver_mux_selector);
			track_1_6_chanY_n11 <= track_1_6_chanY_n11_driver_mux_fanins(track_1_6_chanY_n11_driver_mux_selector);
			track_1_6_chanY_n12 <= track_1_6_chanY_n12_driver_mux_fanins(track_1_6_chanY_n12_driver_mux_selector);
			track_1_6_chanY_n13 <= track_1_6_chanY_n13_driver_mux_fanins(track_1_6_chanY_n13_driver_mux_selector);
			track_1_6_chanY_n14 <= track_1_6_chanY_n14_driver_mux_fanins(track_1_6_chanY_n14_driver_mux_selector);
			track_1_6_chanY_n15 <= track_1_6_chanY_n15_driver_mux_fanins(track_1_6_chanY_n15_driver_mux_selector);
			track_1_6_chanY_n2  <= track_1_6_chanY_n2_driver_mux_fanins(track_1_6_chanY_n2_driver_mux_selector);
			track_1_6_chanY_n3  <= track_1_6_chanY_n3_driver_mux_fanins(track_1_6_chanY_n3_driver_mux_selector);
			track_1_6_chanY_n4  <= track_1_6_chanY_n4_driver_mux_fanins(track_1_6_chanY_n4_driver_mux_selector);
			track_1_6_chanY_n5  <= track_1_6_chanY_n5_driver_mux_fanins(track_1_6_chanY_n5_driver_mux_selector);
			track_1_6_chanY_n6  <= track_1_6_chanY_n6_driver_mux_fanins(track_1_6_chanY_n6_driver_mux_selector);
			track_1_6_chanY_n7  <= track_1_6_chanY_n7_driver_mux_fanins(track_1_6_chanY_n7_driver_mux_selector);
			track_1_6_chanY_n8  <= track_1_6_chanY_n8_driver_mux_fanins(track_1_6_chanY_n8_driver_mux_selector);
			track_1_6_chanY_n9  <= track_1_6_chanY_n9_driver_mux_fanins(track_1_6_chanY_n9_driver_mux_selector);
			track_2_0_chanX_n0  <= track_2_0_chanX_n0_driver_mux_fanins(track_2_0_chanX_n0_driver_mux_selector);
			track_2_0_chanX_n1  <= track_2_0_chanX_n1_driver_mux_fanins(track_2_0_chanX_n1_driver_mux_selector);
			track_2_0_chanX_n10 <= track_2_0_chanX_n10_driver_mux_fanins(track_2_0_chanX_n10_driver_mux_selector);
			track_2_0_chanX_n11 <= track_2_0_chanX_n11_driver_mux_fanins(track_2_0_chanX_n11_driver_mux_selector);
			track_2_0_chanX_n12 <= track_2_0_chanX_n12_driver_mux_fanins(track_2_0_chanX_n12_driver_mux_selector);
			track_2_0_chanX_n13 <= track_2_0_chanX_n13_driver_mux_fanins(track_2_0_chanX_n13_driver_mux_selector);
			track_2_0_chanX_n14 <= track_2_0_chanX_n14_driver_mux_fanins(track_2_0_chanX_n14_driver_mux_selector);
			track_2_0_chanX_n15 <= track_2_0_chanX_n15_driver_mux_fanins(track_2_0_chanX_n15_driver_mux_selector);
			track_2_0_chanX_n2  <= track_2_0_chanX_n2_driver_mux_fanins(track_2_0_chanX_n2_driver_mux_selector);
			track_2_0_chanX_n3  <= track_2_0_chanX_n3_driver_mux_fanins(track_2_0_chanX_n3_driver_mux_selector);
			track_2_0_chanX_n4  <= track_2_0_chanX_n4_driver_mux_fanins(track_2_0_chanX_n4_driver_mux_selector);
			track_2_0_chanX_n5  <= track_2_0_chanX_n5_driver_mux_fanins(track_2_0_chanX_n5_driver_mux_selector);
			track_2_0_chanX_n6  <= track_2_0_chanX_n6_driver_mux_fanins(track_2_0_chanX_n6_driver_mux_selector);
			track_2_0_chanX_n7  <= track_2_0_chanX_n7_driver_mux_fanins(track_2_0_chanX_n7_driver_mux_selector);
			track_2_0_chanX_n8  <= track_2_0_chanX_n8_driver_mux_fanins(track_2_0_chanX_n8_driver_mux_selector);
			track_2_0_chanX_n9  <= track_2_0_chanX_n9_driver_mux_fanins(track_2_0_chanX_n9_driver_mux_selector);
			track_2_1_chanX_n0  <= track_2_1_chanX_n0_driver_mux_fanins(track_2_1_chanX_n0_driver_mux_selector);
			track_2_1_chanX_n1  <= track_2_1_chanX_n1_driver_mux_fanins(track_2_1_chanX_n1_driver_mux_selector);
			track_2_1_chanX_n10 <= track_2_1_chanX_n10_driver_mux_fanins(track_2_1_chanX_n10_driver_mux_selector);
			track_2_1_chanX_n11 <= track_2_1_chanX_n11_driver_mux_fanins(track_2_1_chanX_n11_driver_mux_selector);
			track_2_1_chanX_n12 <= track_2_1_chanX_n12_driver_mux_fanins(track_2_1_chanX_n12_driver_mux_selector);
			track_2_1_chanX_n13 <= track_2_1_chanX_n13_driver_mux_fanins(track_2_1_chanX_n13_driver_mux_selector);
			track_2_1_chanX_n14 <= track_2_1_chanX_n14_driver_mux_fanins(track_2_1_chanX_n14_driver_mux_selector);
			track_2_1_chanX_n15 <= track_2_1_chanX_n15_driver_mux_fanins(track_2_1_chanX_n15_driver_mux_selector);
			track_2_1_chanX_n2  <= track_2_1_chanX_n2_driver_mux_fanins(track_2_1_chanX_n2_driver_mux_selector);
			track_2_1_chanX_n3  <= track_2_1_chanX_n3_driver_mux_fanins(track_2_1_chanX_n3_driver_mux_selector);
			track_2_1_chanX_n4  <= track_2_1_chanX_n4_driver_mux_fanins(track_2_1_chanX_n4_driver_mux_selector);
			track_2_1_chanX_n5  <= track_2_1_chanX_n5_driver_mux_fanins(track_2_1_chanX_n5_driver_mux_selector);
			track_2_1_chanX_n6  <= track_2_1_chanX_n6_driver_mux_fanins(track_2_1_chanX_n6_driver_mux_selector);
			track_2_1_chanX_n7  <= track_2_1_chanX_n7_driver_mux_fanins(track_2_1_chanX_n7_driver_mux_selector);
			track_2_1_chanX_n8  <= track_2_1_chanX_n8_driver_mux_fanins(track_2_1_chanX_n8_driver_mux_selector);
			track_2_1_chanX_n9  <= track_2_1_chanX_n9_driver_mux_fanins(track_2_1_chanX_n9_driver_mux_selector);
			track_2_1_chanY_n0  <= track_2_1_chanY_n0_driver_mux_fanins(track_2_1_chanY_n0_driver_mux_selector);
			track_2_1_chanY_n1  <= track_2_1_chanY_n1_driver_mux_fanins(track_2_1_chanY_n1_driver_mux_selector);
			track_2_1_chanY_n10 <= track_2_1_chanY_n10_driver_mux_fanins(track_2_1_chanY_n10_driver_mux_selector);
			track_2_1_chanY_n11 <= track_2_1_chanY_n11_driver_mux_fanins(track_2_1_chanY_n11_driver_mux_selector);
			track_2_1_chanY_n12 <= track_2_1_chanY_n12_driver_mux_fanins(track_2_1_chanY_n12_driver_mux_selector);
			track_2_1_chanY_n13 <= track_2_1_chanY_n13_driver_mux_fanins(track_2_1_chanY_n13_driver_mux_selector);
			track_2_1_chanY_n14 <= track_2_1_chanY_n14_driver_mux_fanins(track_2_1_chanY_n14_driver_mux_selector);
			track_2_1_chanY_n15 <= track_2_1_chanY_n15_driver_mux_fanins(track_2_1_chanY_n15_driver_mux_selector);
			track_2_1_chanY_n2  <= track_2_1_chanY_n2_driver_mux_fanins(track_2_1_chanY_n2_driver_mux_selector);
			track_2_1_chanY_n3  <= track_2_1_chanY_n3_driver_mux_fanins(track_2_1_chanY_n3_driver_mux_selector);
			track_2_1_chanY_n4  <= track_2_1_chanY_n4_driver_mux_fanins(track_2_1_chanY_n4_driver_mux_selector);
			track_2_1_chanY_n5  <= track_2_1_chanY_n5_driver_mux_fanins(track_2_1_chanY_n5_driver_mux_selector);
			track_2_1_chanY_n6  <= track_2_1_chanY_n6_driver_mux_fanins(track_2_1_chanY_n6_driver_mux_selector);
			track_2_1_chanY_n7  <= track_2_1_chanY_n7_driver_mux_fanins(track_2_1_chanY_n7_driver_mux_selector);
			track_2_1_chanY_n8  <= track_2_1_chanY_n8_driver_mux_fanins(track_2_1_chanY_n8_driver_mux_selector);
			track_2_1_chanY_n9  <= track_2_1_chanY_n9_driver_mux_fanins(track_2_1_chanY_n9_driver_mux_selector);
			track_2_2_chanX_n0  <= track_2_2_chanX_n0_driver_mux_fanins(track_2_2_chanX_n0_driver_mux_selector);
			track_2_2_chanX_n1  <= track_2_2_chanX_n1_driver_mux_fanins(track_2_2_chanX_n1_driver_mux_selector);
			track_2_2_chanX_n10 <= track_2_2_chanX_n10_driver_mux_fanins(track_2_2_chanX_n10_driver_mux_selector);
			track_2_2_chanX_n11 <= track_2_2_chanX_n11_driver_mux_fanins(track_2_2_chanX_n11_driver_mux_selector);
			track_2_2_chanX_n12 <= track_2_2_chanX_n12_driver_mux_fanins(track_2_2_chanX_n12_driver_mux_selector);
			track_2_2_chanX_n13 <= track_2_2_chanX_n13_driver_mux_fanins(track_2_2_chanX_n13_driver_mux_selector);
			track_2_2_chanX_n14 <= track_2_2_chanX_n14_driver_mux_fanins(track_2_2_chanX_n14_driver_mux_selector);
			track_2_2_chanX_n15 <= track_2_2_chanX_n15_driver_mux_fanins(track_2_2_chanX_n15_driver_mux_selector);
			track_2_2_chanX_n2  <= track_2_2_chanX_n2_driver_mux_fanins(track_2_2_chanX_n2_driver_mux_selector);
			track_2_2_chanX_n3  <= track_2_2_chanX_n3_driver_mux_fanins(track_2_2_chanX_n3_driver_mux_selector);
			track_2_2_chanX_n4  <= track_2_2_chanX_n4_driver_mux_fanins(track_2_2_chanX_n4_driver_mux_selector);
			track_2_2_chanX_n5  <= track_2_2_chanX_n5_driver_mux_fanins(track_2_2_chanX_n5_driver_mux_selector);
			track_2_2_chanX_n6  <= track_2_2_chanX_n6_driver_mux_fanins(track_2_2_chanX_n6_driver_mux_selector);
			track_2_2_chanX_n7  <= track_2_2_chanX_n7_driver_mux_fanins(track_2_2_chanX_n7_driver_mux_selector);
			track_2_2_chanX_n8  <= track_2_2_chanX_n8_driver_mux_fanins(track_2_2_chanX_n8_driver_mux_selector);
			track_2_2_chanX_n9  <= track_2_2_chanX_n9_driver_mux_fanins(track_2_2_chanX_n9_driver_mux_selector);
			track_2_2_chanY_n0  <= track_2_2_chanY_n0_driver_mux_fanins(track_2_2_chanY_n0_driver_mux_selector);
			track_2_2_chanY_n1  <= track_2_2_chanY_n1_driver_mux_fanins(track_2_2_chanY_n1_driver_mux_selector);
			track_2_2_chanY_n10 <= track_2_2_chanY_n10_driver_mux_fanins(track_2_2_chanY_n10_driver_mux_selector);
			track_2_2_chanY_n11 <= track_2_2_chanY_n11_driver_mux_fanins(track_2_2_chanY_n11_driver_mux_selector);
			track_2_2_chanY_n12 <= track_2_2_chanY_n12_driver_mux_fanins(track_2_2_chanY_n12_driver_mux_selector);
			track_2_2_chanY_n13 <= track_2_2_chanY_n13_driver_mux_fanins(track_2_2_chanY_n13_driver_mux_selector);
			track_2_2_chanY_n14 <= track_2_2_chanY_n14_driver_mux_fanins(track_2_2_chanY_n14_driver_mux_selector);
			track_2_2_chanY_n15 <= track_2_2_chanY_n15_driver_mux_fanins(track_2_2_chanY_n15_driver_mux_selector);
			track_2_2_chanY_n2  <= track_2_2_chanY_n2_driver_mux_fanins(track_2_2_chanY_n2_driver_mux_selector);
			track_2_2_chanY_n3  <= track_2_2_chanY_n3_driver_mux_fanins(track_2_2_chanY_n3_driver_mux_selector);
			track_2_2_chanY_n4  <= track_2_2_chanY_n4_driver_mux_fanins(track_2_2_chanY_n4_driver_mux_selector);
			track_2_2_chanY_n5  <= track_2_2_chanY_n5_driver_mux_fanins(track_2_2_chanY_n5_driver_mux_selector);
			track_2_2_chanY_n6  <= track_2_2_chanY_n6_driver_mux_fanins(track_2_2_chanY_n6_driver_mux_selector);
			track_2_2_chanY_n7  <= track_2_2_chanY_n7_driver_mux_fanins(track_2_2_chanY_n7_driver_mux_selector);
			track_2_2_chanY_n8  <= track_2_2_chanY_n8_driver_mux_fanins(track_2_2_chanY_n8_driver_mux_selector);
			track_2_2_chanY_n9  <= track_2_2_chanY_n9_driver_mux_fanins(track_2_2_chanY_n9_driver_mux_selector);
			track_2_3_chanX_n0  <= track_2_3_chanX_n0_driver_mux_fanins(track_2_3_chanX_n0_driver_mux_selector);
			track_2_3_chanX_n1  <= track_2_3_chanX_n1_driver_mux_fanins(track_2_3_chanX_n1_driver_mux_selector);
			track_2_3_chanX_n10 <= track_2_3_chanX_n10_driver_mux_fanins(track_2_3_chanX_n10_driver_mux_selector);
			track_2_3_chanX_n11 <= track_2_3_chanX_n11_driver_mux_fanins(track_2_3_chanX_n11_driver_mux_selector);
			track_2_3_chanX_n12 <= track_2_3_chanX_n12_driver_mux_fanins(track_2_3_chanX_n12_driver_mux_selector);
			track_2_3_chanX_n13 <= track_2_3_chanX_n13_driver_mux_fanins(track_2_3_chanX_n13_driver_mux_selector);
			track_2_3_chanX_n14 <= track_2_3_chanX_n14_driver_mux_fanins(track_2_3_chanX_n14_driver_mux_selector);
			track_2_3_chanX_n15 <= track_2_3_chanX_n15_driver_mux_fanins(track_2_3_chanX_n15_driver_mux_selector);
			track_2_3_chanX_n2  <= track_2_3_chanX_n2_driver_mux_fanins(track_2_3_chanX_n2_driver_mux_selector);
			track_2_3_chanX_n3  <= track_2_3_chanX_n3_driver_mux_fanins(track_2_3_chanX_n3_driver_mux_selector);
			track_2_3_chanX_n4  <= track_2_3_chanX_n4_driver_mux_fanins(track_2_3_chanX_n4_driver_mux_selector);
			track_2_3_chanX_n5  <= track_2_3_chanX_n5_driver_mux_fanins(track_2_3_chanX_n5_driver_mux_selector);
			track_2_3_chanX_n6  <= track_2_3_chanX_n6_driver_mux_fanins(track_2_3_chanX_n6_driver_mux_selector);
			track_2_3_chanX_n7  <= track_2_3_chanX_n7_driver_mux_fanins(track_2_3_chanX_n7_driver_mux_selector);
			track_2_3_chanX_n8  <= track_2_3_chanX_n8_driver_mux_fanins(track_2_3_chanX_n8_driver_mux_selector);
			track_2_3_chanX_n9  <= track_2_3_chanX_n9_driver_mux_fanins(track_2_3_chanX_n9_driver_mux_selector);
			track_2_3_chanY_n0  <= track_2_3_chanY_n0_driver_mux_fanins(track_2_3_chanY_n0_driver_mux_selector);
			track_2_3_chanY_n1  <= track_2_3_chanY_n1_driver_mux_fanins(track_2_3_chanY_n1_driver_mux_selector);
			track_2_3_chanY_n10 <= track_2_3_chanY_n10_driver_mux_fanins(track_2_3_chanY_n10_driver_mux_selector);
			track_2_3_chanY_n11 <= track_2_3_chanY_n11_driver_mux_fanins(track_2_3_chanY_n11_driver_mux_selector);
			track_2_3_chanY_n12 <= track_2_3_chanY_n12_driver_mux_fanins(track_2_3_chanY_n12_driver_mux_selector);
			track_2_3_chanY_n13 <= track_2_3_chanY_n13_driver_mux_fanins(track_2_3_chanY_n13_driver_mux_selector);
			track_2_3_chanY_n14 <= track_2_3_chanY_n14_driver_mux_fanins(track_2_3_chanY_n14_driver_mux_selector);
			track_2_3_chanY_n15 <= track_2_3_chanY_n15_driver_mux_fanins(track_2_3_chanY_n15_driver_mux_selector);
			track_2_3_chanY_n2  <= track_2_3_chanY_n2_driver_mux_fanins(track_2_3_chanY_n2_driver_mux_selector);
			track_2_3_chanY_n3  <= track_2_3_chanY_n3_driver_mux_fanins(track_2_3_chanY_n3_driver_mux_selector);
			track_2_3_chanY_n4  <= track_2_3_chanY_n4_driver_mux_fanins(track_2_3_chanY_n4_driver_mux_selector);
			track_2_3_chanY_n5  <= track_2_3_chanY_n5_driver_mux_fanins(track_2_3_chanY_n5_driver_mux_selector);
			track_2_3_chanY_n6  <= track_2_3_chanY_n6_driver_mux_fanins(track_2_3_chanY_n6_driver_mux_selector);
			track_2_3_chanY_n7  <= track_2_3_chanY_n7_driver_mux_fanins(track_2_3_chanY_n7_driver_mux_selector);
			track_2_3_chanY_n8  <= track_2_3_chanY_n8_driver_mux_fanins(track_2_3_chanY_n8_driver_mux_selector);
			track_2_3_chanY_n9  <= track_2_3_chanY_n9_driver_mux_fanins(track_2_3_chanY_n9_driver_mux_selector);
			track_2_4_chanX_n0  <= track_2_4_chanX_n0_driver_mux_fanins(track_2_4_chanX_n0_driver_mux_selector);
			track_2_4_chanX_n1  <= track_2_4_chanX_n1_driver_mux_fanins(track_2_4_chanX_n1_driver_mux_selector);
			track_2_4_chanX_n10 <= track_2_4_chanX_n10_driver_mux_fanins(track_2_4_chanX_n10_driver_mux_selector);
			track_2_4_chanX_n11 <= track_2_4_chanX_n11_driver_mux_fanins(track_2_4_chanX_n11_driver_mux_selector);
			track_2_4_chanX_n12 <= track_2_4_chanX_n12_driver_mux_fanins(track_2_4_chanX_n12_driver_mux_selector);
			track_2_4_chanX_n13 <= track_2_4_chanX_n13_driver_mux_fanins(track_2_4_chanX_n13_driver_mux_selector);
			track_2_4_chanX_n14 <= track_2_4_chanX_n14_driver_mux_fanins(track_2_4_chanX_n14_driver_mux_selector);
			track_2_4_chanX_n15 <= track_2_4_chanX_n15_driver_mux_fanins(track_2_4_chanX_n15_driver_mux_selector);
			track_2_4_chanX_n2  <= track_2_4_chanX_n2_driver_mux_fanins(track_2_4_chanX_n2_driver_mux_selector);
			track_2_4_chanX_n3  <= track_2_4_chanX_n3_driver_mux_fanins(track_2_4_chanX_n3_driver_mux_selector);
			track_2_4_chanX_n4  <= track_2_4_chanX_n4_driver_mux_fanins(track_2_4_chanX_n4_driver_mux_selector);
			track_2_4_chanX_n5  <= track_2_4_chanX_n5_driver_mux_fanins(track_2_4_chanX_n5_driver_mux_selector);
			track_2_4_chanX_n6  <= track_2_4_chanX_n6_driver_mux_fanins(track_2_4_chanX_n6_driver_mux_selector);
			track_2_4_chanX_n7  <= track_2_4_chanX_n7_driver_mux_fanins(track_2_4_chanX_n7_driver_mux_selector);
			track_2_4_chanX_n8  <= track_2_4_chanX_n8_driver_mux_fanins(track_2_4_chanX_n8_driver_mux_selector);
			track_2_4_chanX_n9  <= track_2_4_chanX_n9_driver_mux_fanins(track_2_4_chanX_n9_driver_mux_selector);
			track_2_4_chanY_n0  <= track_2_4_chanY_n0_driver_mux_fanins(track_2_4_chanY_n0_driver_mux_selector);
			track_2_4_chanY_n1  <= track_2_4_chanY_n1_driver_mux_fanins(track_2_4_chanY_n1_driver_mux_selector);
			track_2_4_chanY_n10 <= track_2_4_chanY_n10_driver_mux_fanins(track_2_4_chanY_n10_driver_mux_selector);
			track_2_4_chanY_n11 <= track_2_4_chanY_n11_driver_mux_fanins(track_2_4_chanY_n11_driver_mux_selector);
			track_2_4_chanY_n12 <= track_2_4_chanY_n12_driver_mux_fanins(track_2_4_chanY_n12_driver_mux_selector);
			track_2_4_chanY_n13 <= track_2_4_chanY_n13_driver_mux_fanins(track_2_4_chanY_n13_driver_mux_selector);
			track_2_4_chanY_n14 <= track_2_4_chanY_n14_driver_mux_fanins(track_2_4_chanY_n14_driver_mux_selector);
			track_2_4_chanY_n15 <= track_2_4_chanY_n15_driver_mux_fanins(track_2_4_chanY_n15_driver_mux_selector);
			track_2_4_chanY_n2  <= track_2_4_chanY_n2_driver_mux_fanins(track_2_4_chanY_n2_driver_mux_selector);
			track_2_4_chanY_n3  <= track_2_4_chanY_n3_driver_mux_fanins(track_2_4_chanY_n3_driver_mux_selector);
			track_2_4_chanY_n4  <= track_2_4_chanY_n4_driver_mux_fanins(track_2_4_chanY_n4_driver_mux_selector);
			track_2_4_chanY_n5  <= track_2_4_chanY_n5_driver_mux_fanins(track_2_4_chanY_n5_driver_mux_selector);
			track_2_4_chanY_n6  <= track_2_4_chanY_n6_driver_mux_fanins(track_2_4_chanY_n6_driver_mux_selector);
			track_2_4_chanY_n7  <= track_2_4_chanY_n7_driver_mux_fanins(track_2_4_chanY_n7_driver_mux_selector);
			track_2_4_chanY_n8  <= track_2_4_chanY_n8_driver_mux_fanins(track_2_4_chanY_n8_driver_mux_selector);
			track_2_4_chanY_n9  <= track_2_4_chanY_n9_driver_mux_fanins(track_2_4_chanY_n9_driver_mux_selector);
			track_2_5_chanX_n0  <= track_2_5_chanX_n0_driver_mux_fanins(track_2_5_chanX_n0_driver_mux_selector);
			track_2_5_chanX_n1  <= track_2_5_chanX_n1_driver_mux_fanins(track_2_5_chanX_n1_driver_mux_selector);
			track_2_5_chanX_n10 <= track_2_5_chanX_n10_driver_mux_fanins(track_2_5_chanX_n10_driver_mux_selector);
			track_2_5_chanX_n11 <= track_2_5_chanX_n11_driver_mux_fanins(track_2_5_chanX_n11_driver_mux_selector);
			track_2_5_chanX_n12 <= track_2_5_chanX_n12_driver_mux_fanins(track_2_5_chanX_n12_driver_mux_selector);
			track_2_5_chanX_n13 <= track_2_5_chanX_n13_driver_mux_fanins(track_2_5_chanX_n13_driver_mux_selector);
			track_2_5_chanX_n14 <= track_2_5_chanX_n14_driver_mux_fanins(track_2_5_chanX_n14_driver_mux_selector);
			track_2_5_chanX_n15 <= track_2_5_chanX_n15_driver_mux_fanins(track_2_5_chanX_n15_driver_mux_selector);
			track_2_5_chanX_n2  <= track_2_5_chanX_n2_driver_mux_fanins(track_2_5_chanX_n2_driver_mux_selector);
			track_2_5_chanX_n3  <= track_2_5_chanX_n3_driver_mux_fanins(track_2_5_chanX_n3_driver_mux_selector);
			track_2_5_chanX_n4  <= track_2_5_chanX_n4_driver_mux_fanins(track_2_5_chanX_n4_driver_mux_selector);
			track_2_5_chanX_n5  <= track_2_5_chanX_n5_driver_mux_fanins(track_2_5_chanX_n5_driver_mux_selector);
			track_2_5_chanX_n6  <= track_2_5_chanX_n6_driver_mux_fanins(track_2_5_chanX_n6_driver_mux_selector);
			track_2_5_chanX_n7  <= track_2_5_chanX_n7_driver_mux_fanins(track_2_5_chanX_n7_driver_mux_selector);
			track_2_5_chanX_n8  <= track_2_5_chanX_n8_driver_mux_fanins(track_2_5_chanX_n8_driver_mux_selector);
			track_2_5_chanX_n9  <= track_2_5_chanX_n9_driver_mux_fanins(track_2_5_chanX_n9_driver_mux_selector);
			track_2_5_chanY_n0  <= track_2_5_chanY_n0_driver_mux_fanins(track_2_5_chanY_n0_driver_mux_selector);
			track_2_5_chanY_n1  <= track_2_5_chanY_n1_driver_mux_fanins(track_2_5_chanY_n1_driver_mux_selector);
			track_2_5_chanY_n10 <= track_2_5_chanY_n10_driver_mux_fanins(track_2_5_chanY_n10_driver_mux_selector);
			track_2_5_chanY_n11 <= track_2_5_chanY_n11_driver_mux_fanins(track_2_5_chanY_n11_driver_mux_selector);
			track_2_5_chanY_n12 <= track_2_5_chanY_n12_driver_mux_fanins(track_2_5_chanY_n12_driver_mux_selector);
			track_2_5_chanY_n13 <= track_2_5_chanY_n13_driver_mux_fanins(track_2_5_chanY_n13_driver_mux_selector);
			track_2_5_chanY_n14 <= track_2_5_chanY_n14_driver_mux_fanins(track_2_5_chanY_n14_driver_mux_selector);
			track_2_5_chanY_n15 <= track_2_5_chanY_n15_driver_mux_fanins(track_2_5_chanY_n15_driver_mux_selector);
			track_2_5_chanY_n2  <= track_2_5_chanY_n2_driver_mux_fanins(track_2_5_chanY_n2_driver_mux_selector);
			track_2_5_chanY_n3  <= track_2_5_chanY_n3_driver_mux_fanins(track_2_5_chanY_n3_driver_mux_selector);
			track_2_5_chanY_n4  <= track_2_5_chanY_n4_driver_mux_fanins(track_2_5_chanY_n4_driver_mux_selector);
			track_2_5_chanY_n5  <= track_2_5_chanY_n5_driver_mux_fanins(track_2_5_chanY_n5_driver_mux_selector);
			track_2_5_chanY_n6  <= track_2_5_chanY_n6_driver_mux_fanins(track_2_5_chanY_n6_driver_mux_selector);
			track_2_5_chanY_n7  <= track_2_5_chanY_n7_driver_mux_fanins(track_2_5_chanY_n7_driver_mux_selector);
			track_2_5_chanY_n8  <= track_2_5_chanY_n8_driver_mux_fanins(track_2_5_chanY_n8_driver_mux_selector);
			track_2_5_chanY_n9  <= track_2_5_chanY_n9_driver_mux_fanins(track_2_5_chanY_n9_driver_mux_selector);
			track_2_6_chanX_n0  <= track_2_6_chanX_n0_driver_mux_fanins(track_2_6_chanX_n0_driver_mux_selector);
			track_2_6_chanX_n1  <= track_2_6_chanX_n1_driver_mux_fanins(track_2_6_chanX_n1_driver_mux_selector);
			track_2_6_chanX_n10 <= track_2_6_chanX_n10_driver_mux_fanins(track_2_6_chanX_n10_driver_mux_selector);
			track_2_6_chanX_n11 <= track_2_6_chanX_n11_driver_mux_fanins(track_2_6_chanX_n11_driver_mux_selector);
			track_2_6_chanX_n12 <= track_2_6_chanX_n12_driver_mux_fanins(track_2_6_chanX_n12_driver_mux_selector);
			track_2_6_chanX_n13 <= track_2_6_chanX_n13_driver_mux_fanins(track_2_6_chanX_n13_driver_mux_selector);
			track_2_6_chanX_n14 <= track_2_6_chanX_n14_driver_mux_fanins(track_2_6_chanX_n14_driver_mux_selector);
			track_2_6_chanX_n15 <= track_2_6_chanX_n15_driver_mux_fanins(track_2_6_chanX_n15_driver_mux_selector);
			track_2_6_chanX_n2  <= track_2_6_chanX_n2_driver_mux_fanins(track_2_6_chanX_n2_driver_mux_selector);
			track_2_6_chanX_n3  <= track_2_6_chanX_n3_driver_mux_fanins(track_2_6_chanX_n3_driver_mux_selector);
			track_2_6_chanX_n4  <= track_2_6_chanX_n4_driver_mux_fanins(track_2_6_chanX_n4_driver_mux_selector);
			track_2_6_chanX_n5  <= track_2_6_chanX_n5_driver_mux_fanins(track_2_6_chanX_n5_driver_mux_selector);
			track_2_6_chanX_n6  <= track_2_6_chanX_n6_driver_mux_fanins(track_2_6_chanX_n6_driver_mux_selector);
			track_2_6_chanX_n7  <= track_2_6_chanX_n7_driver_mux_fanins(track_2_6_chanX_n7_driver_mux_selector);
			track_2_6_chanX_n8  <= track_2_6_chanX_n8_driver_mux_fanins(track_2_6_chanX_n8_driver_mux_selector);
			track_2_6_chanX_n9  <= track_2_6_chanX_n9_driver_mux_fanins(track_2_6_chanX_n9_driver_mux_selector);
			track_2_6_chanY_n0  <= track_2_6_chanY_n0_driver_mux_fanins(track_2_6_chanY_n0_driver_mux_selector);
			track_2_6_chanY_n1  <= track_2_6_chanY_n1_driver_mux_fanins(track_2_6_chanY_n1_driver_mux_selector);
			track_2_6_chanY_n10 <= track_2_6_chanY_n10_driver_mux_fanins(track_2_6_chanY_n10_driver_mux_selector);
			track_2_6_chanY_n11 <= track_2_6_chanY_n11_driver_mux_fanins(track_2_6_chanY_n11_driver_mux_selector);
			track_2_6_chanY_n12 <= track_2_6_chanY_n12_driver_mux_fanins(track_2_6_chanY_n12_driver_mux_selector);
			track_2_6_chanY_n13 <= track_2_6_chanY_n13_driver_mux_fanins(track_2_6_chanY_n13_driver_mux_selector);
			track_2_6_chanY_n14 <= track_2_6_chanY_n14_driver_mux_fanins(track_2_6_chanY_n14_driver_mux_selector);
			track_2_6_chanY_n15 <= track_2_6_chanY_n15_driver_mux_fanins(track_2_6_chanY_n15_driver_mux_selector);
			track_2_6_chanY_n2  <= track_2_6_chanY_n2_driver_mux_fanins(track_2_6_chanY_n2_driver_mux_selector);
			track_2_6_chanY_n3  <= track_2_6_chanY_n3_driver_mux_fanins(track_2_6_chanY_n3_driver_mux_selector);
			track_2_6_chanY_n4  <= track_2_6_chanY_n4_driver_mux_fanins(track_2_6_chanY_n4_driver_mux_selector);
			track_2_6_chanY_n5  <= track_2_6_chanY_n5_driver_mux_fanins(track_2_6_chanY_n5_driver_mux_selector);
			track_2_6_chanY_n6  <= track_2_6_chanY_n6_driver_mux_fanins(track_2_6_chanY_n6_driver_mux_selector);
			track_2_6_chanY_n7  <= track_2_6_chanY_n7_driver_mux_fanins(track_2_6_chanY_n7_driver_mux_selector);
			track_2_6_chanY_n8  <= track_2_6_chanY_n8_driver_mux_fanins(track_2_6_chanY_n8_driver_mux_selector);
			track_2_6_chanY_n9  <= track_2_6_chanY_n9_driver_mux_fanins(track_2_6_chanY_n9_driver_mux_selector);
			track_3_0_chanX_n0  <= track_3_0_chanX_n0_driver_mux_fanins(track_3_0_chanX_n0_driver_mux_selector);
			track_3_0_chanX_n1  <= track_3_0_chanX_n1_driver_mux_fanins(track_3_0_chanX_n1_driver_mux_selector);
			track_3_0_chanX_n10 <= track_3_0_chanX_n10_driver_mux_fanins(track_3_0_chanX_n10_driver_mux_selector);
			track_3_0_chanX_n11 <= track_3_0_chanX_n11_driver_mux_fanins(track_3_0_chanX_n11_driver_mux_selector);
			track_3_0_chanX_n12 <= track_3_0_chanX_n12_driver_mux_fanins(track_3_0_chanX_n12_driver_mux_selector);
			track_3_0_chanX_n13 <= track_3_0_chanX_n13_driver_mux_fanins(track_3_0_chanX_n13_driver_mux_selector);
			track_3_0_chanX_n14 <= track_3_0_chanX_n14_driver_mux_fanins(track_3_0_chanX_n14_driver_mux_selector);
			track_3_0_chanX_n15 <= track_3_0_chanX_n15_driver_mux_fanins(track_3_0_chanX_n15_driver_mux_selector);
			track_3_0_chanX_n2  <= track_3_0_chanX_n2_driver_mux_fanins(track_3_0_chanX_n2_driver_mux_selector);
			track_3_0_chanX_n3  <= track_3_0_chanX_n3_driver_mux_fanins(track_3_0_chanX_n3_driver_mux_selector);
			track_3_0_chanX_n4  <= track_3_0_chanX_n4_driver_mux_fanins(track_3_0_chanX_n4_driver_mux_selector);
			track_3_0_chanX_n5  <= track_3_0_chanX_n5_driver_mux_fanins(track_3_0_chanX_n5_driver_mux_selector);
			track_3_0_chanX_n6  <= track_3_0_chanX_n6_driver_mux_fanins(track_3_0_chanX_n6_driver_mux_selector);
			track_3_0_chanX_n7  <= track_3_0_chanX_n7_driver_mux_fanins(track_3_0_chanX_n7_driver_mux_selector);
			track_3_0_chanX_n8  <= track_3_0_chanX_n8_driver_mux_fanins(track_3_0_chanX_n8_driver_mux_selector);
			track_3_0_chanX_n9  <= track_3_0_chanX_n9_driver_mux_fanins(track_3_0_chanX_n9_driver_mux_selector);
			track_3_1_chanX_n0  <= track_3_1_chanX_n0_driver_mux_fanins(track_3_1_chanX_n0_driver_mux_selector);
			track_3_1_chanX_n1  <= track_3_1_chanX_n1_driver_mux_fanins(track_3_1_chanX_n1_driver_mux_selector);
			track_3_1_chanX_n10 <= track_3_1_chanX_n10_driver_mux_fanins(track_3_1_chanX_n10_driver_mux_selector);
			track_3_1_chanX_n11 <= track_3_1_chanX_n11_driver_mux_fanins(track_3_1_chanX_n11_driver_mux_selector);
			track_3_1_chanX_n12 <= track_3_1_chanX_n12_driver_mux_fanins(track_3_1_chanX_n12_driver_mux_selector);
			track_3_1_chanX_n13 <= track_3_1_chanX_n13_driver_mux_fanins(track_3_1_chanX_n13_driver_mux_selector);
			track_3_1_chanX_n14 <= track_3_1_chanX_n14_driver_mux_fanins(track_3_1_chanX_n14_driver_mux_selector);
			track_3_1_chanX_n15 <= track_3_1_chanX_n15_driver_mux_fanins(track_3_1_chanX_n15_driver_mux_selector);
			track_3_1_chanX_n2  <= track_3_1_chanX_n2_driver_mux_fanins(track_3_1_chanX_n2_driver_mux_selector);
			track_3_1_chanX_n3  <= track_3_1_chanX_n3_driver_mux_fanins(track_3_1_chanX_n3_driver_mux_selector);
			track_3_1_chanX_n4  <= track_3_1_chanX_n4_driver_mux_fanins(track_3_1_chanX_n4_driver_mux_selector);
			track_3_1_chanX_n5  <= track_3_1_chanX_n5_driver_mux_fanins(track_3_1_chanX_n5_driver_mux_selector);
			track_3_1_chanX_n6  <= track_3_1_chanX_n6_driver_mux_fanins(track_3_1_chanX_n6_driver_mux_selector);
			track_3_1_chanX_n7  <= track_3_1_chanX_n7_driver_mux_fanins(track_3_1_chanX_n7_driver_mux_selector);
			track_3_1_chanX_n8  <= track_3_1_chanX_n8_driver_mux_fanins(track_3_1_chanX_n8_driver_mux_selector);
			track_3_1_chanX_n9  <= track_3_1_chanX_n9_driver_mux_fanins(track_3_1_chanX_n9_driver_mux_selector);
			track_3_1_chanY_n0  <= track_3_1_chanY_n0_driver_mux_fanins(track_3_1_chanY_n0_driver_mux_selector);
			track_3_1_chanY_n1  <= track_3_1_chanY_n1_driver_mux_fanins(track_3_1_chanY_n1_driver_mux_selector);
			track_3_1_chanY_n10 <= track_3_1_chanY_n10_driver_mux_fanins(track_3_1_chanY_n10_driver_mux_selector);
			track_3_1_chanY_n11 <= track_3_1_chanY_n11_driver_mux_fanins(track_3_1_chanY_n11_driver_mux_selector);
			track_3_1_chanY_n12 <= track_3_1_chanY_n12_driver_mux_fanins(track_3_1_chanY_n12_driver_mux_selector);
			track_3_1_chanY_n13 <= track_3_1_chanY_n13_driver_mux_fanins(track_3_1_chanY_n13_driver_mux_selector);
			track_3_1_chanY_n14 <= track_3_1_chanY_n14_driver_mux_fanins(track_3_1_chanY_n14_driver_mux_selector);
			track_3_1_chanY_n15 <= track_3_1_chanY_n15_driver_mux_fanins(track_3_1_chanY_n15_driver_mux_selector);
			track_3_1_chanY_n2  <= track_3_1_chanY_n2_driver_mux_fanins(track_3_1_chanY_n2_driver_mux_selector);
			track_3_1_chanY_n3  <= track_3_1_chanY_n3_driver_mux_fanins(track_3_1_chanY_n3_driver_mux_selector);
			track_3_1_chanY_n4  <= track_3_1_chanY_n4_driver_mux_fanins(track_3_1_chanY_n4_driver_mux_selector);
			track_3_1_chanY_n5  <= track_3_1_chanY_n5_driver_mux_fanins(track_3_1_chanY_n5_driver_mux_selector);
			track_3_1_chanY_n6  <= track_3_1_chanY_n6_driver_mux_fanins(track_3_1_chanY_n6_driver_mux_selector);
			track_3_1_chanY_n7  <= track_3_1_chanY_n7_driver_mux_fanins(track_3_1_chanY_n7_driver_mux_selector);
			track_3_1_chanY_n8  <= track_3_1_chanY_n8_driver_mux_fanins(track_3_1_chanY_n8_driver_mux_selector);
			track_3_1_chanY_n9  <= track_3_1_chanY_n9_driver_mux_fanins(track_3_1_chanY_n9_driver_mux_selector);
			track_3_2_chanX_n0  <= track_3_2_chanX_n0_driver_mux_fanins(track_3_2_chanX_n0_driver_mux_selector);
			track_3_2_chanX_n1  <= track_3_2_chanX_n1_driver_mux_fanins(track_3_2_chanX_n1_driver_mux_selector);
			track_3_2_chanX_n10 <= track_3_2_chanX_n10_driver_mux_fanins(track_3_2_chanX_n10_driver_mux_selector);
			track_3_2_chanX_n11 <= track_3_2_chanX_n11_driver_mux_fanins(track_3_2_chanX_n11_driver_mux_selector);
			track_3_2_chanX_n12 <= track_3_2_chanX_n12_driver_mux_fanins(track_3_2_chanX_n12_driver_mux_selector);
			track_3_2_chanX_n13 <= track_3_2_chanX_n13_driver_mux_fanins(track_3_2_chanX_n13_driver_mux_selector);
			track_3_2_chanX_n14 <= track_3_2_chanX_n14_driver_mux_fanins(track_3_2_chanX_n14_driver_mux_selector);
			track_3_2_chanX_n15 <= track_3_2_chanX_n15_driver_mux_fanins(track_3_2_chanX_n15_driver_mux_selector);
			track_3_2_chanX_n2  <= track_3_2_chanX_n2_driver_mux_fanins(track_3_2_chanX_n2_driver_mux_selector);
			track_3_2_chanX_n3  <= track_3_2_chanX_n3_driver_mux_fanins(track_3_2_chanX_n3_driver_mux_selector);
			track_3_2_chanX_n4  <= track_3_2_chanX_n4_driver_mux_fanins(track_3_2_chanX_n4_driver_mux_selector);
			track_3_2_chanX_n5  <= track_3_2_chanX_n5_driver_mux_fanins(track_3_2_chanX_n5_driver_mux_selector);
			track_3_2_chanX_n6  <= track_3_2_chanX_n6_driver_mux_fanins(track_3_2_chanX_n6_driver_mux_selector);
			track_3_2_chanX_n7  <= track_3_2_chanX_n7_driver_mux_fanins(track_3_2_chanX_n7_driver_mux_selector);
			track_3_2_chanX_n8  <= track_3_2_chanX_n8_driver_mux_fanins(track_3_2_chanX_n8_driver_mux_selector);
			track_3_2_chanX_n9  <= track_3_2_chanX_n9_driver_mux_fanins(track_3_2_chanX_n9_driver_mux_selector);
			track_3_2_chanY_n0  <= track_3_2_chanY_n0_driver_mux_fanins(track_3_2_chanY_n0_driver_mux_selector);
			track_3_2_chanY_n1  <= track_3_2_chanY_n1_driver_mux_fanins(track_3_2_chanY_n1_driver_mux_selector);
			track_3_2_chanY_n10 <= track_3_2_chanY_n10_driver_mux_fanins(track_3_2_chanY_n10_driver_mux_selector);
			track_3_2_chanY_n11 <= track_3_2_chanY_n11_driver_mux_fanins(track_3_2_chanY_n11_driver_mux_selector);
			track_3_2_chanY_n12 <= track_3_2_chanY_n12_driver_mux_fanins(track_3_2_chanY_n12_driver_mux_selector);
			track_3_2_chanY_n13 <= track_3_2_chanY_n13_driver_mux_fanins(track_3_2_chanY_n13_driver_mux_selector);
			track_3_2_chanY_n14 <= track_3_2_chanY_n14_driver_mux_fanins(track_3_2_chanY_n14_driver_mux_selector);
			track_3_2_chanY_n15 <= track_3_2_chanY_n15_driver_mux_fanins(track_3_2_chanY_n15_driver_mux_selector);
			track_3_2_chanY_n2  <= track_3_2_chanY_n2_driver_mux_fanins(track_3_2_chanY_n2_driver_mux_selector);
			track_3_2_chanY_n3  <= track_3_2_chanY_n3_driver_mux_fanins(track_3_2_chanY_n3_driver_mux_selector);
			track_3_2_chanY_n4  <= track_3_2_chanY_n4_driver_mux_fanins(track_3_2_chanY_n4_driver_mux_selector);
			track_3_2_chanY_n5  <= track_3_2_chanY_n5_driver_mux_fanins(track_3_2_chanY_n5_driver_mux_selector);
			track_3_2_chanY_n6  <= track_3_2_chanY_n6_driver_mux_fanins(track_3_2_chanY_n6_driver_mux_selector);
			track_3_2_chanY_n7  <= track_3_2_chanY_n7_driver_mux_fanins(track_3_2_chanY_n7_driver_mux_selector);
			track_3_2_chanY_n8  <= track_3_2_chanY_n8_driver_mux_fanins(track_3_2_chanY_n8_driver_mux_selector);
			track_3_2_chanY_n9  <= track_3_2_chanY_n9_driver_mux_fanins(track_3_2_chanY_n9_driver_mux_selector);
			track_3_3_chanX_n0  <= track_3_3_chanX_n0_driver_mux_fanins(track_3_3_chanX_n0_driver_mux_selector);
			track_3_3_chanX_n1  <= track_3_3_chanX_n1_driver_mux_fanins(track_3_3_chanX_n1_driver_mux_selector);
			track_3_3_chanX_n10 <= track_3_3_chanX_n10_driver_mux_fanins(track_3_3_chanX_n10_driver_mux_selector);
			track_3_3_chanX_n11 <= track_3_3_chanX_n11_driver_mux_fanins(track_3_3_chanX_n11_driver_mux_selector);
			track_3_3_chanX_n12 <= track_3_3_chanX_n12_driver_mux_fanins(track_3_3_chanX_n12_driver_mux_selector);
			track_3_3_chanX_n13 <= track_3_3_chanX_n13_driver_mux_fanins(track_3_3_chanX_n13_driver_mux_selector);
			track_3_3_chanX_n14 <= track_3_3_chanX_n14_driver_mux_fanins(track_3_3_chanX_n14_driver_mux_selector);
			track_3_3_chanX_n15 <= track_3_3_chanX_n15_driver_mux_fanins(track_3_3_chanX_n15_driver_mux_selector);
			track_3_3_chanX_n2  <= track_3_3_chanX_n2_driver_mux_fanins(track_3_3_chanX_n2_driver_mux_selector);
			track_3_3_chanX_n3  <= track_3_3_chanX_n3_driver_mux_fanins(track_3_3_chanX_n3_driver_mux_selector);
			track_3_3_chanX_n4  <= track_3_3_chanX_n4_driver_mux_fanins(track_3_3_chanX_n4_driver_mux_selector);
			track_3_3_chanX_n5  <= track_3_3_chanX_n5_driver_mux_fanins(track_3_3_chanX_n5_driver_mux_selector);
			track_3_3_chanX_n6  <= track_3_3_chanX_n6_driver_mux_fanins(track_3_3_chanX_n6_driver_mux_selector);
			track_3_3_chanX_n7  <= track_3_3_chanX_n7_driver_mux_fanins(track_3_3_chanX_n7_driver_mux_selector);
			track_3_3_chanX_n8  <= track_3_3_chanX_n8_driver_mux_fanins(track_3_3_chanX_n8_driver_mux_selector);
			track_3_3_chanX_n9  <= track_3_3_chanX_n9_driver_mux_fanins(track_3_3_chanX_n9_driver_mux_selector);
			track_3_3_chanY_n0  <= track_3_3_chanY_n0_driver_mux_fanins(track_3_3_chanY_n0_driver_mux_selector);
			track_3_3_chanY_n1  <= track_3_3_chanY_n1_driver_mux_fanins(track_3_3_chanY_n1_driver_mux_selector);
			track_3_3_chanY_n10 <= track_3_3_chanY_n10_driver_mux_fanins(track_3_3_chanY_n10_driver_mux_selector);
			track_3_3_chanY_n11 <= track_3_3_chanY_n11_driver_mux_fanins(track_3_3_chanY_n11_driver_mux_selector);
			track_3_3_chanY_n12 <= track_3_3_chanY_n12_driver_mux_fanins(track_3_3_chanY_n12_driver_mux_selector);
			track_3_3_chanY_n13 <= track_3_3_chanY_n13_driver_mux_fanins(track_3_3_chanY_n13_driver_mux_selector);
			track_3_3_chanY_n14 <= track_3_3_chanY_n14_driver_mux_fanins(track_3_3_chanY_n14_driver_mux_selector);
			track_3_3_chanY_n15 <= track_3_3_chanY_n15_driver_mux_fanins(track_3_3_chanY_n15_driver_mux_selector);
			track_3_3_chanY_n2  <= track_3_3_chanY_n2_driver_mux_fanins(track_3_3_chanY_n2_driver_mux_selector);
			track_3_3_chanY_n3  <= track_3_3_chanY_n3_driver_mux_fanins(track_3_3_chanY_n3_driver_mux_selector);
			track_3_3_chanY_n4  <= track_3_3_chanY_n4_driver_mux_fanins(track_3_3_chanY_n4_driver_mux_selector);
			track_3_3_chanY_n5  <= track_3_3_chanY_n5_driver_mux_fanins(track_3_3_chanY_n5_driver_mux_selector);
			track_3_3_chanY_n6  <= track_3_3_chanY_n6_driver_mux_fanins(track_3_3_chanY_n6_driver_mux_selector);
			track_3_3_chanY_n7  <= track_3_3_chanY_n7_driver_mux_fanins(track_3_3_chanY_n7_driver_mux_selector);
			track_3_3_chanY_n8  <= track_3_3_chanY_n8_driver_mux_fanins(track_3_3_chanY_n8_driver_mux_selector);
			track_3_3_chanY_n9  <= track_3_3_chanY_n9_driver_mux_fanins(track_3_3_chanY_n9_driver_mux_selector);
			track_3_4_chanX_n0  <= track_3_4_chanX_n0_driver_mux_fanins(track_3_4_chanX_n0_driver_mux_selector);
			track_3_4_chanX_n1  <= track_3_4_chanX_n1_driver_mux_fanins(track_3_4_chanX_n1_driver_mux_selector);
			track_3_4_chanX_n10 <= track_3_4_chanX_n10_driver_mux_fanins(track_3_4_chanX_n10_driver_mux_selector);
			track_3_4_chanX_n11 <= track_3_4_chanX_n11_driver_mux_fanins(track_3_4_chanX_n11_driver_mux_selector);
			track_3_4_chanX_n12 <= track_3_4_chanX_n12_driver_mux_fanins(track_3_4_chanX_n12_driver_mux_selector);
			track_3_4_chanX_n13 <= track_3_4_chanX_n13_driver_mux_fanins(track_3_4_chanX_n13_driver_mux_selector);
			track_3_4_chanX_n14 <= track_3_4_chanX_n14_driver_mux_fanins(track_3_4_chanX_n14_driver_mux_selector);
			track_3_4_chanX_n15 <= track_3_4_chanX_n15_driver_mux_fanins(track_3_4_chanX_n15_driver_mux_selector);
			track_3_4_chanX_n2  <= track_3_4_chanX_n2_driver_mux_fanins(track_3_4_chanX_n2_driver_mux_selector);
			track_3_4_chanX_n3  <= track_3_4_chanX_n3_driver_mux_fanins(track_3_4_chanX_n3_driver_mux_selector);
			track_3_4_chanX_n4  <= track_3_4_chanX_n4_driver_mux_fanins(track_3_4_chanX_n4_driver_mux_selector);
			track_3_4_chanX_n5  <= track_3_4_chanX_n5_driver_mux_fanins(track_3_4_chanX_n5_driver_mux_selector);
			track_3_4_chanX_n6  <= track_3_4_chanX_n6_driver_mux_fanins(track_3_4_chanX_n6_driver_mux_selector);
			track_3_4_chanX_n7  <= track_3_4_chanX_n7_driver_mux_fanins(track_3_4_chanX_n7_driver_mux_selector);
			track_3_4_chanX_n8  <= track_3_4_chanX_n8_driver_mux_fanins(track_3_4_chanX_n8_driver_mux_selector);
			track_3_4_chanX_n9  <= track_3_4_chanX_n9_driver_mux_fanins(track_3_4_chanX_n9_driver_mux_selector);
			track_3_4_chanY_n0  <= track_3_4_chanY_n0_driver_mux_fanins(track_3_4_chanY_n0_driver_mux_selector);
			track_3_4_chanY_n1  <= track_3_4_chanY_n1_driver_mux_fanins(track_3_4_chanY_n1_driver_mux_selector);
			track_3_4_chanY_n10 <= track_3_4_chanY_n10_driver_mux_fanins(track_3_4_chanY_n10_driver_mux_selector);
			track_3_4_chanY_n11 <= track_3_4_chanY_n11_driver_mux_fanins(track_3_4_chanY_n11_driver_mux_selector);
			track_3_4_chanY_n12 <= track_3_4_chanY_n12_driver_mux_fanins(track_3_4_chanY_n12_driver_mux_selector);
			track_3_4_chanY_n13 <= track_3_4_chanY_n13_driver_mux_fanins(track_3_4_chanY_n13_driver_mux_selector);
			track_3_4_chanY_n14 <= track_3_4_chanY_n14_driver_mux_fanins(track_3_4_chanY_n14_driver_mux_selector);
			track_3_4_chanY_n15 <= track_3_4_chanY_n15_driver_mux_fanins(track_3_4_chanY_n15_driver_mux_selector);
			track_3_4_chanY_n2  <= track_3_4_chanY_n2_driver_mux_fanins(track_3_4_chanY_n2_driver_mux_selector);
			track_3_4_chanY_n3  <= track_3_4_chanY_n3_driver_mux_fanins(track_3_4_chanY_n3_driver_mux_selector);
			track_3_4_chanY_n4  <= track_3_4_chanY_n4_driver_mux_fanins(track_3_4_chanY_n4_driver_mux_selector);
			track_3_4_chanY_n5  <= track_3_4_chanY_n5_driver_mux_fanins(track_3_4_chanY_n5_driver_mux_selector);
			track_3_4_chanY_n6  <= track_3_4_chanY_n6_driver_mux_fanins(track_3_4_chanY_n6_driver_mux_selector);
			track_3_4_chanY_n7  <= track_3_4_chanY_n7_driver_mux_fanins(track_3_4_chanY_n7_driver_mux_selector);
			track_3_4_chanY_n8  <= track_3_4_chanY_n8_driver_mux_fanins(track_3_4_chanY_n8_driver_mux_selector);
			track_3_4_chanY_n9  <= track_3_4_chanY_n9_driver_mux_fanins(track_3_4_chanY_n9_driver_mux_selector);
			track_3_5_chanX_n0  <= track_3_5_chanX_n0_driver_mux_fanins(track_3_5_chanX_n0_driver_mux_selector);
			track_3_5_chanX_n1  <= track_3_5_chanX_n1_driver_mux_fanins(track_3_5_chanX_n1_driver_mux_selector);
			track_3_5_chanX_n10 <= track_3_5_chanX_n10_driver_mux_fanins(track_3_5_chanX_n10_driver_mux_selector);
			track_3_5_chanX_n11 <= track_3_5_chanX_n11_driver_mux_fanins(track_3_5_chanX_n11_driver_mux_selector);
			track_3_5_chanX_n12 <= track_3_5_chanX_n12_driver_mux_fanins(track_3_5_chanX_n12_driver_mux_selector);
			track_3_5_chanX_n13 <= track_3_5_chanX_n13_driver_mux_fanins(track_3_5_chanX_n13_driver_mux_selector);
			track_3_5_chanX_n14 <= track_3_5_chanX_n14_driver_mux_fanins(track_3_5_chanX_n14_driver_mux_selector);
			track_3_5_chanX_n15 <= track_3_5_chanX_n15_driver_mux_fanins(track_3_5_chanX_n15_driver_mux_selector);
			track_3_5_chanX_n2  <= track_3_5_chanX_n2_driver_mux_fanins(track_3_5_chanX_n2_driver_mux_selector);
			track_3_5_chanX_n3  <= track_3_5_chanX_n3_driver_mux_fanins(track_3_5_chanX_n3_driver_mux_selector);
			track_3_5_chanX_n4  <= track_3_5_chanX_n4_driver_mux_fanins(track_3_5_chanX_n4_driver_mux_selector);
			track_3_5_chanX_n5  <= track_3_5_chanX_n5_driver_mux_fanins(track_3_5_chanX_n5_driver_mux_selector);
			track_3_5_chanX_n6  <= track_3_5_chanX_n6_driver_mux_fanins(track_3_5_chanX_n6_driver_mux_selector);
			track_3_5_chanX_n7  <= track_3_5_chanX_n7_driver_mux_fanins(track_3_5_chanX_n7_driver_mux_selector);
			track_3_5_chanX_n8  <= track_3_5_chanX_n8_driver_mux_fanins(track_3_5_chanX_n8_driver_mux_selector);
			track_3_5_chanX_n9  <= track_3_5_chanX_n9_driver_mux_fanins(track_3_5_chanX_n9_driver_mux_selector);
			track_3_5_chanY_n0  <= track_3_5_chanY_n0_driver_mux_fanins(track_3_5_chanY_n0_driver_mux_selector);
			track_3_5_chanY_n1  <= track_3_5_chanY_n1_driver_mux_fanins(track_3_5_chanY_n1_driver_mux_selector);
			track_3_5_chanY_n10 <= track_3_5_chanY_n10_driver_mux_fanins(track_3_5_chanY_n10_driver_mux_selector);
			track_3_5_chanY_n11 <= track_3_5_chanY_n11_driver_mux_fanins(track_3_5_chanY_n11_driver_mux_selector);
			track_3_5_chanY_n12 <= track_3_5_chanY_n12_driver_mux_fanins(track_3_5_chanY_n12_driver_mux_selector);
			track_3_5_chanY_n13 <= track_3_5_chanY_n13_driver_mux_fanins(track_3_5_chanY_n13_driver_mux_selector);
			track_3_5_chanY_n14 <= track_3_5_chanY_n14_driver_mux_fanins(track_3_5_chanY_n14_driver_mux_selector);
			track_3_5_chanY_n15 <= track_3_5_chanY_n15_driver_mux_fanins(track_3_5_chanY_n15_driver_mux_selector);
			track_3_5_chanY_n2  <= track_3_5_chanY_n2_driver_mux_fanins(track_3_5_chanY_n2_driver_mux_selector);
			track_3_5_chanY_n3  <= track_3_5_chanY_n3_driver_mux_fanins(track_3_5_chanY_n3_driver_mux_selector);
			track_3_5_chanY_n4  <= track_3_5_chanY_n4_driver_mux_fanins(track_3_5_chanY_n4_driver_mux_selector);
			track_3_5_chanY_n5  <= track_3_5_chanY_n5_driver_mux_fanins(track_3_5_chanY_n5_driver_mux_selector);
			track_3_5_chanY_n6  <= track_3_5_chanY_n6_driver_mux_fanins(track_3_5_chanY_n6_driver_mux_selector);
			track_3_5_chanY_n7  <= track_3_5_chanY_n7_driver_mux_fanins(track_3_5_chanY_n7_driver_mux_selector);
			track_3_5_chanY_n8  <= track_3_5_chanY_n8_driver_mux_fanins(track_3_5_chanY_n8_driver_mux_selector);
			track_3_5_chanY_n9  <= track_3_5_chanY_n9_driver_mux_fanins(track_3_5_chanY_n9_driver_mux_selector);
			track_3_6_chanX_n0  <= track_3_6_chanX_n0_driver_mux_fanins(track_3_6_chanX_n0_driver_mux_selector);
			track_3_6_chanX_n1  <= track_3_6_chanX_n1_driver_mux_fanins(track_3_6_chanX_n1_driver_mux_selector);
			track_3_6_chanX_n10 <= track_3_6_chanX_n10_driver_mux_fanins(track_3_6_chanX_n10_driver_mux_selector);
			track_3_6_chanX_n11 <= track_3_6_chanX_n11_driver_mux_fanins(track_3_6_chanX_n11_driver_mux_selector);
			track_3_6_chanX_n12 <= track_3_6_chanX_n12_driver_mux_fanins(track_3_6_chanX_n12_driver_mux_selector);
			track_3_6_chanX_n13 <= track_3_6_chanX_n13_driver_mux_fanins(track_3_6_chanX_n13_driver_mux_selector);
			track_3_6_chanX_n14 <= track_3_6_chanX_n14_driver_mux_fanins(track_3_6_chanX_n14_driver_mux_selector);
			track_3_6_chanX_n15 <= track_3_6_chanX_n15_driver_mux_fanins(track_3_6_chanX_n15_driver_mux_selector);
			track_3_6_chanX_n2  <= track_3_6_chanX_n2_driver_mux_fanins(track_3_6_chanX_n2_driver_mux_selector);
			track_3_6_chanX_n3  <= track_3_6_chanX_n3_driver_mux_fanins(track_3_6_chanX_n3_driver_mux_selector);
			track_3_6_chanX_n4  <= track_3_6_chanX_n4_driver_mux_fanins(track_3_6_chanX_n4_driver_mux_selector);
			track_3_6_chanX_n5  <= track_3_6_chanX_n5_driver_mux_fanins(track_3_6_chanX_n5_driver_mux_selector);
			track_3_6_chanX_n6  <= track_3_6_chanX_n6_driver_mux_fanins(track_3_6_chanX_n6_driver_mux_selector);
			track_3_6_chanX_n7  <= track_3_6_chanX_n7_driver_mux_fanins(track_3_6_chanX_n7_driver_mux_selector);
			track_3_6_chanX_n8  <= track_3_6_chanX_n8_driver_mux_fanins(track_3_6_chanX_n8_driver_mux_selector);
			track_3_6_chanX_n9  <= track_3_6_chanX_n9_driver_mux_fanins(track_3_6_chanX_n9_driver_mux_selector);
			track_3_6_chanY_n0  <= track_3_6_chanY_n0_driver_mux_fanins(track_3_6_chanY_n0_driver_mux_selector);
			track_3_6_chanY_n1  <= track_3_6_chanY_n1_driver_mux_fanins(track_3_6_chanY_n1_driver_mux_selector);
			track_3_6_chanY_n10 <= track_3_6_chanY_n10_driver_mux_fanins(track_3_6_chanY_n10_driver_mux_selector);
			track_3_6_chanY_n11 <= track_3_6_chanY_n11_driver_mux_fanins(track_3_6_chanY_n11_driver_mux_selector);
			track_3_6_chanY_n12 <= track_3_6_chanY_n12_driver_mux_fanins(track_3_6_chanY_n12_driver_mux_selector);
			track_3_6_chanY_n13 <= track_3_6_chanY_n13_driver_mux_fanins(track_3_6_chanY_n13_driver_mux_selector);
			track_3_6_chanY_n14 <= track_3_6_chanY_n14_driver_mux_fanins(track_3_6_chanY_n14_driver_mux_selector);
			track_3_6_chanY_n15 <= track_3_6_chanY_n15_driver_mux_fanins(track_3_6_chanY_n15_driver_mux_selector);
			track_3_6_chanY_n2  <= track_3_6_chanY_n2_driver_mux_fanins(track_3_6_chanY_n2_driver_mux_selector);
			track_3_6_chanY_n3  <= track_3_6_chanY_n3_driver_mux_fanins(track_3_6_chanY_n3_driver_mux_selector);
			track_3_6_chanY_n4  <= track_3_6_chanY_n4_driver_mux_fanins(track_3_6_chanY_n4_driver_mux_selector);
			track_3_6_chanY_n5  <= track_3_6_chanY_n5_driver_mux_fanins(track_3_6_chanY_n5_driver_mux_selector);
			track_3_6_chanY_n6  <= track_3_6_chanY_n6_driver_mux_fanins(track_3_6_chanY_n6_driver_mux_selector);
			track_3_6_chanY_n7  <= track_3_6_chanY_n7_driver_mux_fanins(track_3_6_chanY_n7_driver_mux_selector);
			track_3_6_chanY_n8  <= track_3_6_chanY_n8_driver_mux_fanins(track_3_6_chanY_n8_driver_mux_selector);
			track_3_6_chanY_n9  <= track_3_6_chanY_n9_driver_mux_fanins(track_3_6_chanY_n9_driver_mux_selector);
			track_4_0_chanX_n0  <= track_4_0_chanX_n0_driver_mux_fanins(track_4_0_chanX_n0_driver_mux_selector);
			track_4_0_chanX_n1  <= track_4_0_chanX_n1_driver_mux_fanins(track_4_0_chanX_n1_driver_mux_selector);
			track_4_0_chanX_n10 <= track_4_0_chanX_n10_driver_mux_fanins(track_4_0_chanX_n10_driver_mux_selector);
			track_4_0_chanX_n11 <= track_4_0_chanX_n11_driver_mux_fanins(track_4_0_chanX_n11_driver_mux_selector);
			track_4_0_chanX_n12 <= track_4_0_chanX_n12_driver_mux_fanins(track_4_0_chanX_n12_driver_mux_selector);
			track_4_0_chanX_n13 <= track_4_0_chanX_n13_driver_mux_fanins(track_4_0_chanX_n13_driver_mux_selector);
			track_4_0_chanX_n14 <= track_4_0_chanX_n14_driver_mux_fanins(track_4_0_chanX_n14_driver_mux_selector);
			track_4_0_chanX_n15 <= track_4_0_chanX_n15_driver_mux_fanins(track_4_0_chanX_n15_driver_mux_selector);
			track_4_0_chanX_n2  <= track_4_0_chanX_n2_driver_mux_fanins(track_4_0_chanX_n2_driver_mux_selector);
			track_4_0_chanX_n3  <= track_4_0_chanX_n3_driver_mux_fanins(track_4_0_chanX_n3_driver_mux_selector);
			track_4_0_chanX_n4  <= track_4_0_chanX_n4_driver_mux_fanins(track_4_0_chanX_n4_driver_mux_selector);
			track_4_0_chanX_n5  <= track_4_0_chanX_n5_driver_mux_fanins(track_4_0_chanX_n5_driver_mux_selector);
			track_4_0_chanX_n6  <= track_4_0_chanX_n6_driver_mux_fanins(track_4_0_chanX_n6_driver_mux_selector);
			track_4_0_chanX_n7  <= track_4_0_chanX_n7_driver_mux_fanins(track_4_0_chanX_n7_driver_mux_selector);
			track_4_0_chanX_n8  <= track_4_0_chanX_n8_driver_mux_fanins(track_4_0_chanX_n8_driver_mux_selector);
			track_4_0_chanX_n9  <= track_4_0_chanX_n9_driver_mux_fanins(track_4_0_chanX_n9_driver_mux_selector);
			track_4_1_chanX_n0  <= track_4_1_chanX_n0_driver_mux_fanins(track_4_1_chanX_n0_driver_mux_selector);
			track_4_1_chanX_n1  <= track_4_1_chanX_n1_driver_mux_fanins(track_4_1_chanX_n1_driver_mux_selector);
			track_4_1_chanX_n10 <= track_4_1_chanX_n10_driver_mux_fanins(track_4_1_chanX_n10_driver_mux_selector);
			track_4_1_chanX_n11 <= track_4_1_chanX_n11_driver_mux_fanins(track_4_1_chanX_n11_driver_mux_selector);
			track_4_1_chanX_n12 <= track_4_1_chanX_n12_driver_mux_fanins(track_4_1_chanX_n12_driver_mux_selector);
			track_4_1_chanX_n13 <= track_4_1_chanX_n13_driver_mux_fanins(track_4_1_chanX_n13_driver_mux_selector);
			track_4_1_chanX_n14 <= track_4_1_chanX_n14_driver_mux_fanins(track_4_1_chanX_n14_driver_mux_selector);
			track_4_1_chanX_n15 <= track_4_1_chanX_n15_driver_mux_fanins(track_4_1_chanX_n15_driver_mux_selector);
			track_4_1_chanX_n2  <= track_4_1_chanX_n2_driver_mux_fanins(track_4_1_chanX_n2_driver_mux_selector);
			track_4_1_chanX_n3  <= track_4_1_chanX_n3_driver_mux_fanins(track_4_1_chanX_n3_driver_mux_selector);
			track_4_1_chanX_n4  <= track_4_1_chanX_n4_driver_mux_fanins(track_4_1_chanX_n4_driver_mux_selector);
			track_4_1_chanX_n5  <= track_4_1_chanX_n5_driver_mux_fanins(track_4_1_chanX_n5_driver_mux_selector);
			track_4_1_chanX_n6  <= track_4_1_chanX_n6_driver_mux_fanins(track_4_1_chanX_n6_driver_mux_selector);
			track_4_1_chanX_n7  <= track_4_1_chanX_n7_driver_mux_fanins(track_4_1_chanX_n7_driver_mux_selector);
			track_4_1_chanX_n8  <= track_4_1_chanX_n8_driver_mux_fanins(track_4_1_chanX_n8_driver_mux_selector);
			track_4_1_chanX_n9  <= track_4_1_chanX_n9_driver_mux_fanins(track_4_1_chanX_n9_driver_mux_selector);
			track_4_1_chanY_n0  <= track_4_1_chanY_n0_driver_mux_fanins(track_4_1_chanY_n0_driver_mux_selector);
			track_4_1_chanY_n1  <= track_4_1_chanY_n1_driver_mux_fanins(track_4_1_chanY_n1_driver_mux_selector);
			track_4_1_chanY_n10 <= track_4_1_chanY_n10_driver_mux_fanins(track_4_1_chanY_n10_driver_mux_selector);
			track_4_1_chanY_n11 <= track_4_1_chanY_n11_driver_mux_fanins(track_4_1_chanY_n11_driver_mux_selector);
			track_4_1_chanY_n12 <= track_4_1_chanY_n12_driver_mux_fanins(track_4_1_chanY_n12_driver_mux_selector);
			track_4_1_chanY_n13 <= track_4_1_chanY_n13_driver_mux_fanins(track_4_1_chanY_n13_driver_mux_selector);
			track_4_1_chanY_n14 <= track_4_1_chanY_n14_driver_mux_fanins(track_4_1_chanY_n14_driver_mux_selector);
			track_4_1_chanY_n15 <= track_4_1_chanY_n15_driver_mux_fanins(track_4_1_chanY_n15_driver_mux_selector);
			track_4_1_chanY_n2  <= track_4_1_chanY_n2_driver_mux_fanins(track_4_1_chanY_n2_driver_mux_selector);
			track_4_1_chanY_n3  <= track_4_1_chanY_n3_driver_mux_fanins(track_4_1_chanY_n3_driver_mux_selector);
			track_4_1_chanY_n4  <= track_4_1_chanY_n4_driver_mux_fanins(track_4_1_chanY_n4_driver_mux_selector);
			track_4_1_chanY_n5  <= track_4_1_chanY_n5_driver_mux_fanins(track_4_1_chanY_n5_driver_mux_selector);
			track_4_1_chanY_n6  <= track_4_1_chanY_n6_driver_mux_fanins(track_4_1_chanY_n6_driver_mux_selector);
			track_4_1_chanY_n7  <= track_4_1_chanY_n7_driver_mux_fanins(track_4_1_chanY_n7_driver_mux_selector);
			track_4_1_chanY_n8  <= track_4_1_chanY_n8_driver_mux_fanins(track_4_1_chanY_n8_driver_mux_selector);
			track_4_1_chanY_n9  <= track_4_1_chanY_n9_driver_mux_fanins(track_4_1_chanY_n9_driver_mux_selector);
			track_4_2_chanX_n0  <= track_4_2_chanX_n0_driver_mux_fanins(track_4_2_chanX_n0_driver_mux_selector);
			track_4_2_chanX_n1  <= track_4_2_chanX_n1_driver_mux_fanins(track_4_2_chanX_n1_driver_mux_selector);
			track_4_2_chanX_n10 <= track_4_2_chanX_n10_driver_mux_fanins(track_4_2_chanX_n10_driver_mux_selector);
			track_4_2_chanX_n11 <= track_4_2_chanX_n11_driver_mux_fanins(track_4_2_chanX_n11_driver_mux_selector);
			track_4_2_chanX_n12 <= track_4_2_chanX_n12_driver_mux_fanins(track_4_2_chanX_n12_driver_mux_selector);
			track_4_2_chanX_n13 <= track_4_2_chanX_n13_driver_mux_fanins(track_4_2_chanX_n13_driver_mux_selector);
			track_4_2_chanX_n14 <= track_4_2_chanX_n14_driver_mux_fanins(track_4_2_chanX_n14_driver_mux_selector);
			track_4_2_chanX_n15 <= track_4_2_chanX_n15_driver_mux_fanins(track_4_2_chanX_n15_driver_mux_selector);
			track_4_2_chanX_n2  <= track_4_2_chanX_n2_driver_mux_fanins(track_4_2_chanX_n2_driver_mux_selector);
			track_4_2_chanX_n3  <= track_4_2_chanX_n3_driver_mux_fanins(track_4_2_chanX_n3_driver_mux_selector);
			track_4_2_chanX_n4  <= track_4_2_chanX_n4_driver_mux_fanins(track_4_2_chanX_n4_driver_mux_selector);
			track_4_2_chanX_n5  <= track_4_2_chanX_n5_driver_mux_fanins(track_4_2_chanX_n5_driver_mux_selector);
			track_4_2_chanX_n6  <= track_4_2_chanX_n6_driver_mux_fanins(track_4_2_chanX_n6_driver_mux_selector);
			track_4_2_chanX_n7  <= track_4_2_chanX_n7_driver_mux_fanins(track_4_2_chanX_n7_driver_mux_selector);
			track_4_2_chanX_n8  <= track_4_2_chanX_n8_driver_mux_fanins(track_4_2_chanX_n8_driver_mux_selector);
			track_4_2_chanX_n9  <= track_4_2_chanX_n9_driver_mux_fanins(track_4_2_chanX_n9_driver_mux_selector);
			track_4_2_chanY_n0  <= track_4_2_chanY_n0_driver_mux_fanins(track_4_2_chanY_n0_driver_mux_selector);
			track_4_2_chanY_n1  <= track_4_2_chanY_n1_driver_mux_fanins(track_4_2_chanY_n1_driver_mux_selector);
			track_4_2_chanY_n10 <= track_4_2_chanY_n10_driver_mux_fanins(track_4_2_chanY_n10_driver_mux_selector);
			track_4_2_chanY_n11 <= track_4_2_chanY_n11_driver_mux_fanins(track_4_2_chanY_n11_driver_mux_selector);
			track_4_2_chanY_n12 <= track_4_2_chanY_n12_driver_mux_fanins(track_4_2_chanY_n12_driver_mux_selector);
			track_4_2_chanY_n13 <= track_4_2_chanY_n13_driver_mux_fanins(track_4_2_chanY_n13_driver_mux_selector);
			track_4_2_chanY_n14 <= track_4_2_chanY_n14_driver_mux_fanins(track_4_2_chanY_n14_driver_mux_selector);
			track_4_2_chanY_n15 <= track_4_2_chanY_n15_driver_mux_fanins(track_4_2_chanY_n15_driver_mux_selector);
			track_4_2_chanY_n2  <= track_4_2_chanY_n2_driver_mux_fanins(track_4_2_chanY_n2_driver_mux_selector);
			track_4_2_chanY_n3  <= track_4_2_chanY_n3_driver_mux_fanins(track_4_2_chanY_n3_driver_mux_selector);
			track_4_2_chanY_n4  <= track_4_2_chanY_n4_driver_mux_fanins(track_4_2_chanY_n4_driver_mux_selector);
			track_4_2_chanY_n5  <= track_4_2_chanY_n5_driver_mux_fanins(track_4_2_chanY_n5_driver_mux_selector);
			track_4_2_chanY_n6  <= track_4_2_chanY_n6_driver_mux_fanins(track_4_2_chanY_n6_driver_mux_selector);
			track_4_2_chanY_n7  <= track_4_2_chanY_n7_driver_mux_fanins(track_4_2_chanY_n7_driver_mux_selector);
			track_4_2_chanY_n8  <= track_4_2_chanY_n8_driver_mux_fanins(track_4_2_chanY_n8_driver_mux_selector);
			track_4_2_chanY_n9  <= track_4_2_chanY_n9_driver_mux_fanins(track_4_2_chanY_n9_driver_mux_selector);
			track_4_3_chanX_n0  <= track_4_3_chanX_n0_driver_mux_fanins(track_4_3_chanX_n0_driver_mux_selector);
			track_4_3_chanX_n1  <= track_4_3_chanX_n1_driver_mux_fanins(track_4_3_chanX_n1_driver_mux_selector);
			track_4_3_chanX_n10 <= track_4_3_chanX_n10_driver_mux_fanins(track_4_3_chanX_n10_driver_mux_selector);
			track_4_3_chanX_n11 <= track_4_3_chanX_n11_driver_mux_fanins(track_4_3_chanX_n11_driver_mux_selector);
			track_4_3_chanX_n12 <= track_4_3_chanX_n12_driver_mux_fanins(track_4_3_chanX_n12_driver_mux_selector);
			track_4_3_chanX_n13 <= track_4_3_chanX_n13_driver_mux_fanins(track_4_3_chanX_n13_driver_mux_selector);
			track_4_3_chanX_n14 <= track_4_3_chanX_n14_driver_mux_fanins(track_4_3_chanX_n14_driver_mux_selector);
			track_4_3_chanX_n15 <= track_4_3_chanX_n15_driver_mux_fanins(track_4_3_chanX_n15_driver_mux_selector);
			track_4_3_chanX_n2  <= track_4_3_chanX_n2_driver_mux_fanins(track_4_3_chanX_n2_driver_mux_selector);
			track_4_3_chanX_n3  <= track_4_3_chanX_n3_driver_mux_fanins(track_4_3_chanX_n3_driver_mux_selector);
			track_4_3_chanX_n4  <= track_4_3_chanX_n4_driver_mux_fanins(track_4_3_chanX_n4_driver_mux_selector);
			track_4_3_chanX_n5  <= track_4_3_chanX_n5_driver_mux_fanins(track_4_3_chanX_n5_driver_mux_selector);
			track_4_3_chanX_n6  <= track_4_3_chanX_n6_driver_mux_fanins(track_4_3_chanX_n6_driver_mux_selector);
			track_4_3_chanX_n7  <= track_4_3_chanX_n7_driver_mux_fanins(track_4_3_chanX_n7_driver_mux_selector);
			track_4_3_chanX_n8  <= track_4_3_chanX_n8_driver_mux_fanins(track_4_3_chanX_n8_driver_mux_selector);
			track_4_3_chanX_n9  <= track_4_3_chanX_n9_driver_mux_fanins(track_4_3_chanX_n9_driver_mux_selector);
			track_4_3_chanY_n0  <= track_4_3_chanY_n0_driver_mux_fanins(track_4_3_chanY_n0_driver_mux_selector);
			track_4_3_chanY_n1  <= track_4_3_chanY_n1_driver_mux_fanins(track_4_3_chanY_n1_driver_mux_selector);
			track_4_3_chanY_n10 <= track_4_3_chanY_n10_driver_mux_fanins(track_4_3_chanY_n10_driver_mux_selector);
			track_4_3_chanY_n11 <= track_4_3_chanY_n11_driver_mux_fanins(track_4_3_chanY_n11_driver_mux_selector);
			track_4_3_chanY_n12 <= track_4_3_chanY_n12_driver_mux_fanins(track_4_3_chanY_n12_driver_mux_selector);
			track_4_3_chanY_n13 <= track_4_3_chanY_n13_driver_mux_fanins(track_4_3_chanY_n13_driver_mux_selector);
			track_4_3_chanY_n14 <= track_4_3_chanY_n14_driver_mux_fanins(track_4_3_chanY_n14_driver_mux_selector);
			track_4_3_chanY_n15 <= track_4_3_chanY_n15_driver_mux_fanins(track_4_3_chanY_n15_driver_mux_selector);
			track_4_3_chanY_n2  <= track_4_3_chanY_n2_driver_mux_fanins(track_4_3_chanY_n2_driver_mux_selector);
			track_4_3_chanY_n3  <= track_4_3_chanY_n3_driver_mux_fanins(track_4_3_chanY_n3_driver_mux_selector);
			track_4_3_chanY_n4  <= track_4_3_chanY_n4_driver_mux_fanins(track_4_3_chanY_n4_driver_mux_selector);
			track_4_3_chanY_n5  <= track_4_3_chanY_n5_driver_mux_fanins(track_4_3_chanY_n5_driver_mux_selector);
			track_4_3_chanY_n6  <= track_4_3_chanY_n6_driver_mux_fanins(track_4_3_chanY_n6_driver_mux_selector);
			track_4_3_chanY_n7  <= track_4_3_chanY_n7_driver_mux_fanins(track_4_3_chanY_n7_driver_mux_selector);
			track_4_3_chanY_n8  <= track_4_3_chanY_n8_driver_mux_fanins(track_4_3_chanY_n8_driver_mux_selector);
			track_4_3_chanY_n9  <= track_4_3_chanY_n9_driver_mux_fanins(track_4_3_chanY_n9_driver_mux_selector);
			track_4_4_chanX_n0  <= track_4_4_chanX_n0_driver_mux_fanins(track_4_4_chanX_n0_driver_mux_selector);
			track_4_4_chanX_n1  <= track_4_4_chanX_n1_driver_mux_fanins(track_4_4_chanX_n1_driver_mux_selector);
			track_4_4_chanX_n10 <= track_4_4_chanX_n10_driver_mux_fanins(track_4_4_chanX_n10_driver_mux_selector);
			track_4_4_chanX_n11 <= track_4_4_chanX_n11_driver_mux_fanins(track_4_4_chanX_n11_driver_mux_selector);
			track_4_4_chanX_n12 <= track_4_4_chanX_n12_driver_mux_fanins(track_4_4_chanX_n12_driver_mux_selector);
			track_4_4_chanX_n13 <= track_4_4_chanX_n13_driver_mux_fanins(track_4_4_chanX_n13_driver_mux_selector);
			track_4_4_chanX_n14 <= track_4_4_chanX_n14_driver_mux_fanins(track_4_4_chanX_n14_driver_mux_selector);
			track_4_4_chanX_n15 <= track_4_4_chanX_n15_driver_mux_fanins(track_4_4_chanX_n15_driver_mux_selector);
			track_4_4_chanX_n2  <= track_4_4_chanX_n2_driver_mux_fanins(track_4_4_chanX_n2_driver_mux_selector);
			track_4_4_chanX_n3  <= track_4_4_chanX_n3_driver_mux_fanins(track_4_4_chanX_n3_driver_mux_selector);
			track_4_4_chanX_n4  <= track_4_4_chanX_n4_driver_mux_fanins(track_4_4_chanX_n4_driver_mux_selector);
			track_4_4_chanX_n5  <= track_4_4_chanX_n5_driver_mux_fanins(track_4_4_chanX_n5_driver_mux_selector);
			track_4_4_chanX_n6  <= track_4_4_chanX_n6_driver_mux_fanins(track_4_4_chanX_n6_driver_mux_selector);
			track_4_4_chanX_n7  <= track_4_4_chanX_n7_driver_mux_fanins(track_4_4_chanX_n7_driver_mux_selector);
			track_4_4_chanX_n8  <= track_4_4_chanX_n8_driver_mux_fanins(track_4_4_chanX_n8_driver_mux_selector);
			track_4_4_chanX_n9  <= track_4_4_chanX_n9_driver_mux_fanins(track_4_4_chanX_n9_driver_mux_selector);
			track_4_4_chanY_n0  <= track_4_4_chanY_n0_driver_mux_fanins(track_4_4_chanY_n0_driver_mux_selector);
			track_4_4_chanY_n1  <= track_4_4_chanY_n1_driver_mux_fanins(track_4_4_chanY_n1_driver_mux_selector);
			track_4_4_chanY_n10 <= track_4_4_chanY_n10_driver_mux_fanins(track_4_4_chanY_n10_driver_mux_selector);
			track_4_4_chanY_n11 <= track_4_4_chanY_n11_driver_mux_fanins(track_4_4_chanY_n11_driver_mux_selector);
			track_4_4_chanY_n12 <= track_4_4_chanY_n12_driver_mux_fanins(track_4_4_chanY_n12_driver_mux_selector);
			track_4_4_chanY_n13 <= track_4_4_chanY_n13_driver_mux_fanins(track_4_4_chanY_n13_driver_mux_selector);
			track_4_4_chanY_n14 <= track_4_4_chanY_n14_driver_mux_fanins(track_4_4_chanY_n14_driver_mux_selector);
			track_4_4_chanY_n15 <= track_4_4_chanY_n15_driver_mux_fanins(track_4_4_chanY_n15_driver_mux_selector);
			track_4_4_chanY_n2  <= track_4_4_chanY_n2_driver_mux_fanins(track_4_4_chanY_n2_driver_mux_selector);
			track_4_4_chanY_n3  <= track_4_4_chanY_n3_driver_mux_fanins(track_4_4_chanY_n3_driver_mux_selector);
			track_4_4_chanY_n4  <= track_4_4_chanY_n4_driver_mux_fanins(track_4_4_chanY_n4_driver_mux_selector);
			track_4_4_chanY_n5  <= track_4_4_chanY_n5_driver_mux_fanins(track_4_4_chanY_n5_driver_mux_selector);
			track_4_4_chanY_n6  <= track_4_4_chanY_n6_driver_mux_fanins(track_4_4_chanY_n6_driver_mux_selector);
			track_4_4_chanY_n7  <= track_4_4_chanY_n7_driver_mux_fanins(track_4_4_chanY_n7_driver_mux_selector);
			track_4_4_chanY_n8  <= track_4_4_chanY_n8_driver_mux_fanins(track_4_4_chanY_n8_driver_mux_selector);
			track_4_4_chanY_n9  <= track_4_4_chanY_n9_driver_mux_fanins(track_4_4_chanY_n9_driver_mux_selector);
			track_4_5_chanX_n0  <= track_4_5_chanX_n0_driver_mux_fanins(track_4_5_chanX_n0_driver_mux_selector);
			track_4_5_chanX_n1  <= track_4_5_chanX_n1_driver_mux_fanins(track_4_5_chanX_n1_driver_mux_selector);
			track_4_5_chanX_n10 <= track_4_5_chanX_n10_driver_mux_fanins(track_4_5_chanX_n10_driver_mux_selector);
			track_4_5_chanX_n11 <= track_4_5_chanX_n11_driver_mux_fanins(track_4_5_chanX_n11_driver_mux_selector);
			track_4_5_chanX_n12 <= track_4_5_chanX_n12_driver_mux_fanins(track_4_5_chanX_n12_driver_mux_selector);
			track_4_5_chanX_n13 <= track_4_5_chanX_n13_driver_mux_fanins(track_4_5_chanX_n13_driver_mux_selector);
			track_4_5_chanX_n14 <= track_4_5_chanX_n14_driver_mux_fanins(track_4_5_chanX_n14_driver_mux_selector);
			track_4_5_chanX_n15 <= track_4_5_chanX_n15_driver_mux_fanins(track_4_5_chanX_n15_driver_mux_selector);
			track_4_5_chanX_n2  <= track_4_5_chanX_n2_driver_mux_fanins(track_4_5_chanX_n2_driver_mux_selector);
			track_4_5_chanX_n3  <= track_4_5_chanX_n3_driver_mux_fanins(track_4_5_chanX_n3_driver_mux_selector);
			track_4_5_chanX_n4  <= track_4_5_chanX_n4_driver_mux_fanins(track_4_5_chanX_n4_driver_mux_selector);
			track_4_5_chanX_n5  <= track_4_5_chanX_n5_driver_mux_fanins(track_4_5_chanX_n5_driver_mux_selector);
			track_4_5_chanX_n6  <= track_4_5_chanX_n6_driver_mux_fanins(track_4_5_chanX_n6_driver_mux_selector);
			track_4_5_chanX_n7  <= track_4_5_chanX_n7_driver_mux_fanins(track_4_5_chanX_n7_driver_mux_selector);
			track_4_5_chanX_n8  <= track_4_5_chanX_n8_driver_mux_fanins(track_4_5_chanX_n8_driver_mux_selector);
			track_4_5_chanX_n9  <= track_4_5_chanX_n9_driver_mux_fanins(track_4_5_chanX_n9_driver_mux_selector);
			track_4_5_chanY_n0  <= track_4_5_chanY_n0_driver_mux_fanins(track_4_5_chanY_n0_driver_mux_selector);
			track_4_5_chanY_n1  <= track_4_5_chanY_n1_driver_mux_fanins(track_4_5_chanY_n1_driver_mux_selector);
			track_4_5_chanY_n10 <= track_4_5_chanY_n10_driver_mux_fanins(track_4_5_chanY_n10_driver_mux_selector);
			track_4_5_chanY_n11 <= track_4_5_chanY_n11_driver_mux_fanins(track_4_5_chanY_n11_driver_mux_selector);
			track_4_5_chanY_n12 <= track_4_5_chanY_n12_driver_mux_fanins(track_4_5_chanY_n12_driver_mux_selector);
			track_4_5_chanY_n13 <= track_4_5_chanY_n13_driver_mux_fanins(track_4_5_chanY_n13_driver_mux_selector);
			track_4_5_chanY_n14 <= track_4_5_chanY_n14_driver_mux_fanins(track_4_5_chanY_n14_driver_mux_selector);
			track_4_5_chanY_n15 <= track_4_5_chanY_n15_driver_mux_fanins(track_4_5_chanY_n15_driver_mux_selector);
			track_4_5_chanY_n2  <= track_4_5_chanY_n2_driver_mux_fanins(track_4_5_chanY_n2_driver_mux_selector);
			track_4_5_chanY_n3  <= track_4_5_chanY_n3_driver_mux_fanins(track_4_5_chanY_n3_driver_mux_selector);
			track_4_5_chanY_n4  <= track_4_5_chanY_n4_driver_mux_fanins(track_4_5_chanY_n4_driver_mux_selector);
			track_4_5_chanY_n5  <= track_4_5_chanY_n5_driver_mux_fanins(track_4_5_chanY_n5_driver_mux_selector);
			track_4_5_chanY_n6  <= track_4_5_chanY_n6_driver_mux_fanins(track_4_5_chanY_n6_driver_mux_selector);
			track_4_5_chanY_n7  <= track_4_5_chanY_n7_driver_mux_fanins(track_4_5_chanY_n7_driver_mux_selector);
			track_4_5_chanY_n8  <= track_4_5_chanY_n8_driver_mux_fanins(track_4_5_chanY_n8_driver_mux_selector);
			track_4_5_chanY_n9  <= track_4_5_chanY_n9_driver_mux_fanins(track_4_5_chanY_n9_driver_mux_selector);
			track_4_6_chanX_n0  <= track_4_6_chanX_n0_driver_mux_fanins(track_4_6_chanX_n0_driver_mux_selector);
			track_4_6_chanX_n1  <= track_4_6_chanX_n1_driver_mux_fanins(track_4_6_chanX_n1_driver_mux_selector);
			track_4_6_chanX_n10 <= track_4_6_chanX_n10_driver_mux_fanins(track_4_6_chanX_n10_driver_mux_selector);
			track_4_6_chanX_n11 <= track_4_6_chanX_n11_driver_mux_fanins(track_4_6_chanX_n11_driver_mux_selector);
			track_4_6_chanX_n12 <= track_4_6_chanX_n12_driver_mux_fanins(track_4_6_chanX_n12_driver_mux_selector);
			track_4_6_chanX_n13 <= track_4_6_chanX_n13_driver_mux_fanins(track_4_6_chanX_n13_driver_mux_selector);
			track_4_6_chanX_n14 <= track_4_6_chanX_n14_driver_mux_fanins(track_4_6_chanX_n14_driver_mux_selector);
			track_4_6_chanX_n15 <= track_4_6_chanX_n15_driver_mux_fanins(track_4_6_chanX_n15_driver_mux_selector);
			track_4_6_chanX_n2  <= track_4_6_chanX_n2_driver_mux_fanins(track_4_6_chanX_n2_driver_mux_selector);
			track_4_6_chanX_n3  <= track_4_6_chanX_n3_driver_mux_fanins(track_4_6_chanX_n3_driver_mux_selector);
			track_4_6_chanX_n4  <= track_4_6_chanX_n4_driver_mux_fanins(track_4_6_chanX_n4_driver_mux_selector);
			track_4_6_chanX_n5  <= track_4_6_chanX_n5_driver_mux_fanins(track_4_6_chanX_n5_driver_mux_selector);
			track_4_6_chanX_n6  <= track_4_6_chanX_n6_driver_mux_fanins(track_4_6_chanX_n6_driver_mux_selector);
			track_4_6_chanX_n7  <= track_4_6_chanX_n7_driver_mux_fanins(track_4_6_chanX_n7_driver_mux_selector);
			track_4_6_chanX_n8  <= track_4_6_chanX_n8_driver_mux_fanins(track_4_6_chanX_n8_driver_mux_selector);
			track_4_6_chanX_n9  <= track_4_6_chanX_n9_driver_mux_fanins(track_4_6_chanX_n9_driver_mux_selector);
			track_4_6_chanY_n0  <= track_4_6_chanY_n0_driver_mux_fanins(track_4_6_chanY_n0_driver_mux_selector);
			track_4_6_chanY_n1  <= track_4_6_chanY_n1_driver_mux_fanins(track_4_6_chanY_n1_driver_mux_selector);
			track_4_6_chanY_n10 <= track_4_6_chanY_n10_driver_mux_fanins(track_4_6_chanY_n10_driver_mux_selector);
			track_4_6_chanY_n11 <= track_4_6_chanY_n11_driver_mux_fanins(track_4_6_chanY_n11_driver_mux_selector);
			track_4_6_chanY_n12 <= track_4_6_chanY_n12_driver_mux_fanins(track_4_6_chanY_n12_driver_mux_selector);
			track_4_6_chanY_n13 <= track_4_6_chanY_n13_driver_mux_fanins(track_4_6_chanY_n13_driver_mux_selector);
			track_4_6_chanY_n14 <= track_4_6_chanY_n14_driver_mux_fanins(track_4_6_chanY_n14_driver_mux_selector);
			track_4_6_chanY_n15 <= track_4_6_chanY_n15_driver_mux_fanins(track_4_6_chanY_n15_driver_mux_selector);
			track_4_6_chanY_n2  <= track_4_6_chanY_n2_driver_mux_fanins(track_4_6_chanY_n2_driver_mux_selector);
			track_4_6_chanY_n3  <= track_4_6_chanY_n3_driver_mux_fanins(track_4_6_chanY_n3_driver_mux_selector);
			track_4_6_chanY_n4  <= track_4_6_chanY_n4_driver_mux_fanins(track_4_6_chanY_n4_driver_mux_selector);
			track_4_6_chanY_n5  <= track_4_6_chanY_n5_driver_mux_fanins(track_4_6_chanY_n5_driver_mux_selector);
			track_4_6_chanY_n6  <= track_4_6_chanY_n6_driver_mux_fanins(track_4_6_chanY_n6_driver_mux_selector);
			track_4_6_chanY_n7  <= track_4_6_chanY_n7_driver_mux_fanins(track_4_6_chanY_n7_driver_mux_selector);
			track_4_6_chanY_n8  <= track_4_6_chanY_n8_driver_mux_fanins(track_4_6_chanY_n8_driver_mux_selector);
			track_4_6_chanY_n9  <= track_4_6_chanY_n9_driver_mux_fanins(track_4_6_chanY_n9_driver_mux_selector);
			track_5_0_chanX_n0  <= track_5_0_chanX_n0_driver_mux_fanins(track_5_0_chanX_n0_driver_mux_selector);
			track_5_0_chanX_n1  <= track_5_0_chanX_n1_driver_mux_fanins(track_5_0_chanX_n1_driver_mux_selector);
			track_5_0_chanX_n10 <= track_5_0_chanX_n10_driver_mux_fanins(track_5_0_chanX_n10_driver_mux_selector);
			track_5_0_chanX_n11 <= track_5_0_chanX_n11_driver_mux_fanins(track_5_0_chanX_n11_driver_mux_selector);
			track_5_0_chanX_n12 <= track_5_0_chanX_n12_driver_mux_fanins(track_5_0_chanX_n12_driver_mux_selector);
			track_5_0_chanX_n13 <= track_5_0_chanX_n13_driver_mux_fanins(track_5_0_chanX_n13_driver_mux_selector);
			track_5_0_chanX_n14 <= track_5_0_chanX_n14_driver_mux_fanins(track_5_0_chanX_n14_driver_mux_selector);
			track_5_0_chanX_n15 <= track_5_0_chanX_n15_driver_mux_fanins(track_5_0_chanX_n15_driver_mux_selector);
			track_5_0_chanX_n2  <= track_5_0_chanX_n2_driver_mux_fanins(track_5_0_chanX_n2_driver_mux_selector);
			track_5_0_chanX_n3  <= track_5_0_chanX_n3_driver_mux_fanins(track_5_0_chanX_n3_driver_mux_selector);
			track_5_0_chanX_n4  <= track_5_0_chanX_n4_driver_mux_fanins(track_5_0_chanX_n4_driver_mux_selector);
			track_5_0_chanX_n5  <= track_5_0_chanX_n5_driver_mux_fanins(track_5_0_chanX_n5_driver_mux_selector);
			track_5_0_chanX_n6  <= track_5_0_chanX_n6_driver_mux_fanins(track_5_0_chanX_n6_driver_mux_selector);
			track_5_0_chanX_n7  <= track_5_0_chanX_n7_driver_mux_fanins(track_5_0_chanX_n7_driver_mux_selector);
			track_5_0_chanX_n8  <= track_5_0_chanX_n8_driver_mux_fanins(track_5_0_chanX_n8_driver_mux_selector);
			track_5_0_chanX_n9  <= track_5_0_chanX_n9_driver_mux_fanins(track_5_0_chanX_n9_driver_mux_selector);
			track_5_1_chanX_n0  <= track_5_1_chanX_n0_driver_mux_fanins(track_5_1_chanX_n0_driver_mux_selector);
			track_5_1_chanX_n1  <= track_5_1_chanX_n1_driver_mux_fanins(track_5_1_chanX_n1_driver_mux_selector);
			track_5_1_chanX_n10 <= track_5_1_chanX_n10_driver_mux_fanins(track_5_1_chanX_n10_driver_mux_selector);
			track_5_1_chanX_n11 <= track_5_1_chanX_n11_driver_mux_fanins(track_5_1_chanX_n11_driver_mux_selector);
			track_5_1_chanX_n12 <= track_5_1_chanX_n12_driver_mux_fanins(track_5_1_chanX_n12_driver_mux_selector);
			track_5_1_chanX_n13 <= track_5_1_chanX_n13_driver_mux_fanins(track_5_1_chanX_n13_driver_mux_selector);
			track_5_1_chanX_n14 <= track_5_1_chanX_n14_driver_mux_fanins(track_5_1_chanX_n14_driver_mux_selector);
			track_5_1_chanX_n15 <= track_5_1_chanX_n15_driver_mux_fanins(track_5_1_chanX_n15_driver_mux_selector);
			track_5_1_chanX_n2  <= track_5_1_chanX_n2_driver_mux_fanins(track_5_1_chanX_n2_driver_mux_selector);
			track_5_1_chanX_n3  <= track_5_1_chanX_n3_driver_mux_fanins(track_5_1_chanX_n3_driver_mux_selector);
			track_5_1_chanX_n4  <= track_5_1_chanX_n4_driver_mux_fanins(track_5_1_chanX_n4_driver_mux_selector);
			track_5_1_chanX_n5  <= track_5_1_chanX_n5_driver_mux_fanins(track_5_1_chanX_n5_driver_mux_selector);
			track_5_1_chanX_n6  <= track_5_1_chanX_n6_driver_mux_fanins(track_5_1_chanX_n6_driver_mux_selector);
			track_5_1_chanX_n7  <= track_5_1_chanX_n7_driver_mux_fanins(track_5_1_chanX_n7_driver_mux_selector);
			track_5_1_chanX_n8  <= track_5_1_chanX_n8_driver_mux_fanins(track_5_1_chanX_n8_driver_mux_selector);
			track_5_1_chanX_n9  <= track_5_1_chanX_n9_driver_mux_fanins(track_5_1_chanX_n9_driver_mux_selector);
			track_5_1_chanY_n0  <= track_5_1_chanY_n0_driver_mux_fanins(track_5_1_chanY_n0_driver_mux_selector);
			track_5_1_chanY_n1  <= track_5_1_chanY_n1_driver_mux_fanins(track_5_1_chanY_n1_driver_mux_selector);
			track_5_1_chanY_n10 <= track_5_1_chanY_n10_driver_mux_fanins(track_5_1_chanY_n10_driver_mux_selector);
			track_5_1_chanY_n11 <= track_5_1_chanY_n11_driver_mux_fanins(track_5_1_chanY_n11_driver_mux_selector);
			track_5_1_chanY_n12 <= track_5_1_chanY_n12_driver_mux_fanins(track_5_1_chanY_n12_driver_mux_selector);
			track_5_1_chanY_n13 <= track_5_1_chanY_n13_driver_mux_fanins(track_5_1_chanY_n13_driver_mux_selector);
			track_5_1_chanY_n14 <= track_5_1_chanY_n14_driver_mux_fanins(track_5_1_chanY_n14_driver_mux_selector);
			track_5_1_chanY_n15 <= track_5_1_chanY_n15_driver_mux_fanins(track_5_1_chanY_n15_driver_mux_selector);
			track_5_1_chanY_n2  <= track_5_1_chanY_n2_driver_mux_fanins(track_5_1_chanY_n2_driver_mux_selector);
			track_5_1_chanY_n3  <= track_5_1_chanY_n3_driver_mux_fanins(track_5_1_chanY_n3_driver_mux_selector);
			track_5_1_chanY_n4  <= track_5_1_chanY_n4_driver_mux_fanins(track_5_1_chanY_n4_driver_mux_selector);
			track_5_1_chanY_n5  <= track_5_1_chanY_n5_driver_mux_fanins(track_5_1_chanY_n5_driver_mux_selector);
			track_5_1_chanY_n6  <= track_5_1_chanY_n6_driver_mux_fanins(track_5_1_chanY_n6_driver_mux_selector);
			track_5_1_chanY_n7  <= track_5_1_chanY_n7_driver_mux_fanins(track_5_1_chanY_n7_driver_mux_selector);
			track_5_1_chanY_n8  <= track_5_1_chanY_n8_driver_mux_fanins(track_5_1_chanY_n8_driver_mux_selector);
			track_5_1_chanY_n9  <= track_5_1_chanY_n9_driver_mux_fanins(track_5_1_chanY_n9_driver_mux_selector);
			track_5_2_chanX_n0  <= track_5_2_chanX_n0_driver_mux_fanins(track_5_2_chanX_n0_driver_mux_selector);
			track_5_2_chanX_n1  <= track_5_2_chanX_n1_driver_mux_fanins(track_5_2_chanX_n1_driver_mux_selector);
			track_5_2_chanX_n10 <= track_5_2_chanX_n10_driver_mux_fanins(track_5_2_chanX_n10_driver_mux_selector);
			track_5_2_chanX_n11 <= track_5_2_chanX_n11_driver_mux_fanins(track_5_2_chanX_n11_driver_mux_selector);
			track_5_2_chanX_n12 <= track_5_2_chanX_n12_driver_mux_fanins(track_5_2_chanX_n12_driver_mux_selector);
			track_5_2_chanX_n13 <= track_5_2_chanX_n13_driver_mux_fanins(track_5_2_chanX_n13_driver_mux_selector);
			track_5_2_chanX_n14 <= track_5_2_chanX_n14_driver_mux_fanins(track_5_2_chanX_n14_driver_mux_selector);
			track_5_2_chanX_n15 <= track_5_2_chanX_n15_driver_mux_fanins(track_5_2_chanX_n15_driver_mux_selector);
			track_5_2_chanX_n2  <= track_5_2_chanX_n2_driver_mux_fanins(track_5_2_chanX_n2_driver_mux_selector);
			track_5_2_chanX_n3  <= track_5_2_chanX_n3_driver_mux_fanins(track_5_2_chanX_n3_driver_mux_selector);
			track_5_2_chanX_n4  <= track_5_2_chanX_n4_driver_mux_fanins(track_5_2_chanX_n4_driver_mux_selector);
			track_5_2_chanX_n5  <= track_5_2_chanX_n5_driver_mux_fanins(track_5_2_chanX_n5_driver_mux_selector);
			track_5_2_chanX_n6  <= track_5_2_chanX_n6_driver_mux_fanins(track_5_2_chanX_n6_driver_mux_selector);
			track_5_2_chanX_n7  <= track_5_2_chanX_n7_driver_mux_fanins(track_5_2_chanX_n7_driver_mux_selector);
			track_5_2_chanX_n8  <= track_5_2_chanX_n8_driver_mux_fanins(track_5_2_chanX_n8_driver_mux_selector);
			track_5_2_chanX_n9  <= track_5_2_chanX_n9_driver_mux_fanins(track_5_2_chanX_n9_driver_mux_selector);
			track_5_2_chanY_n0  <= track_5_2_chanY_n0_driver_mux_fanins(track_5_2_chanY_n0_driver_mux_selector);
			track_5_2_chanY_n1  <= track_5_2_chanY_n1_driver_mux_fanins(track_5_2_chanY_n1_driver_mux_selector);
			track_5_2_chanY_n10 <= track_5_2_chanY_n10_driver_mux_fanins(track_5_2_chanY_n10_driver_mux_selector);
			track_5_2_chanY_n11 <= track_5_2_chanY_n11_driver_mux_fanins(track_5_2_chanY_n11_driver_mux_selector);
			track_5_2_chanY_n12 <= track_5_2_chanY_n12_driver_mux_fanins(track_5_2_chanY_n12_driver_mux_selector);
			track_5_2_chanY_n13 <= track_5_2_chanY_n13_driver_mux_fanins(track_5_2_chanY_n13_driver_mux_selector);
			track_5_2_chanY_n14 <= track_5_2_chanY_n14_driver_mux_fanins(track_5_2_chanY_n14_driver_mux_selector);
			track_5_2_chanY_n15 <= track_5_2_chanY_n15_driver_mux_fanins(track_5_2_chanY_n15_driver_mux_selector);
			track_5_2_chanY_n2  <= track_5_2_chanY_n2_driver_mux_fanins(track_5_2_chanY_n2_driver_mux_selector);
			track_5_2_chanY_n3  <= track_5_2_chanY_n3_driver_mux_fanins(track_5_2_chanY_n3_driver_mux_selector);
			track_5_2_chanY_n4  <= track_5_2_chanY_n4_driver_mux_fanins(track_5_2_chanY_n4_driver_mux_selector);
			track_5_2_chanY_n5  <= track_5_2_chanY_n5_driver_mux_fanins(track_5_2_chanY_n5_driver_mux_selector);
			track_5_2_chanY_n6  <= track_5_2_chanY_n6_driver_mux_fanins(track_5_2_chanY_n6_driver_mux_selector);
			track_5_2_chanY_n7  <= track_5_2_chanY_n7_driver_mux_fanins(track_5_2_chanY_n7_driver_mux_selector);
			track_5_2_chanY_n8  <= track_5_2_chanY_n8_driver_mux_fanins(track_5_2_chanY_n8_driver_mux_selector);
			track_5_2_chanY_n9  <= track_5_2_chanY_n9_driver_mux_fanins(track_5_2_chanY_n9_driver_mux_selector);
			track_5_3_chanX_n0  <= track_5_3_chanX_n0_driver_mux_fanins(track_5_3_chanX_n0_driver_mux_selector);
			track_5_3_chanX_n1  <= track_5_3_chanX_n1_driver_mux_fanins(track_5_3_chanX_n1_driver_mux_selector);
			track_5_3_chanX_n10 <= track_5_3_chanX_n10_driver_mux_fanins(track_5_3_chanX_n10_driver_mux_selector);
			track_5_3_chanX_n11 <= track_5_3_chanX_n11_driver_mux_fanins(track_5_3_chanX_n11_driver_mux_selector);
			track_5_3_chanX_n12 <= track_5_3_chanX_n12_driver_mux_fanins(track_5_3_chanX_n12_driver_mux_selector);
			track_5_3_chanX_n13 <= track_5_3_chanX_n13_driver_mux_fanins(track_5_3_chanX_n13_driver_mux_selector);
			track_5_3_chanX_n14 <= track_5_3_chanX_n14_driver_mux_fanins(track_5_3_chanX_n14_driver_mux_selector);
			track_5_3_chanX_n15 <= track_5_3_chanX_n15_driver_mux_fanins(track_5_3_chanX_n15_driver_mux_selector);
			track_5_3_chanX_n2  <= track_5_3_chanX_n2_driver_mux_fanins(track_5_3_chanX_n2_driver_mux_selector);
			track_5_3_chanX_n3  <= track_5_3_chanX_n3_driver_mux_fanins(track_5_3_chanX_n3_driver_mux_selector);
			track_5_3_chanX_n4  <= track_5_3_chanX_n4_driver_mux_fanins(track_5_3_chanX_n4_driver_mux_selector);
			track_5_3_chanX_n5  <= track_5_3_chanX_n5_driver_mux_fanins(track_5_3_chanX_n5_driver_mux_selector);
			track_5_3_chanX_n6  <= track_5_3_chanX_n6_driver_mux_fanins(track_5_3_chanX_n6_driver_mux_selector);
			track_5_3_chanX_n7  <= track_5_3_chanX_n7_driver_mux_fanins(track_5_3_chanX_n7_driver_mux_selector);
			track_5_3_chanX_n8  <= track_5_3_chanX_n8_driver_mux_fanins(track_5_3_chanX_n8_driver_mux_selector);
			track_5_3_chanX_n9  <= track_5_3_chanX_n9_driver_mux_fanins(track_5_3_chanX_n9_driver_mux_selector);
			track_5_3_chanY_n0  <= track_5_3_chanY_n0_driver_mux_fanins(track_5_3_chanY_n0_driver_mux_selector);
			track_5_3_chanY_n1  <= track_5_3_chanY_n1_driver_mux_fanins(track_5_3_chanY_n1_driver_mux_selector);
			track_5_3_chanY_n10 <= track_5_3_chanY_n10_driver_mux_fanins(track_5_3_chanY_n10_driver_mux_selector);
			track_5_3_chanY_n11 <= track_5_3_chanY_n11_driver_mux_fanins(track_5_3_chanY_n11_driver_mux_selector);
			track_5_3_chanY_n12 <= track_5_3_chanY_n12_driver_mux_fanins(track_5_3_chanY_n12_driver_mux_selector);
			track_5_3_chanY_n13 <= track_5_3_chanY_n13_driver_mux_fanins(track_5_3_chanY_n13_driver_mux_selector);
			track_5_3_chanY_n14 <= track_5_3_chanY_n14_driver_mux_fanins(track_5_3_chanY_n14_driver_mux_selector);
			track_5_3_chanY_n15 <= track_5_3_chanY_n15_driver_mux_fanins(track_5_3_chanY_n15_driver_mux_selector);
			track_5_3_chanY_n2  <= track_5_3_chanY_n2_driver_mux_fanins(track_5_3_chanY_n2_driver_mux_selector);
			track_5_3_chanY_n3  <= track_5_3_chanY_n3_driver_mux_fanins(track_5_3_chanY_n3_driver_mux_selector);
			track_5_3_chanY_n4  <= track_5_3_chanY_n4_driver_mux_fanins(track_5_3_chanY_n4_driver_mux_selector);
			track_5_3_chanY_n5  <= track_5_3_chanY_n5_driver_mux_fanins(track_5_3_chanY_n5_driver_mux_selector);
			track_5_3_chanY_n6  <= track_5_3_chanY_n6_driver_mux_fanins(track_5_3_chanY_n6_driver_mux_selector);
			track_5_3_chanY_n7  <= track_5_3_chanY_n7_driver_mux_fanins(track_5_3_chanY_n7_driver_mux_selector);
			track_5_3_chanY_n8  <= track_5_3_chanY_n8_driver_mux_fanins(track_5_3_chanY_n8_driver_mux_selector);
			track_5_3_chanY_n9  <= track_5_3_chanY_n9_driver_mux_fanins(track_5_3_chanY_n9_driver_mux_selector);
			track_5_4_chanX_n0  <= track_5_4_chanX_n0_driver_mux_fanins(track_5_4_chanX_n0_driver_mux_selector);
			track_5_4_chanX_n1  <= track_5_4_chanX_n1_driver_mux_fanins(track_5_4_chanX_n1_driver_mux_selector);
			track_5_4_chanX_n10 <= track_5_4_chanX_n10_driver_mux_fanins(track_5_4_chanX_n10_driver_mux_selector);
			track_5_4_chanX_n11 <= track_5_4_chanX_n11_driver_mux_fanins(track_5_4_chanX_n11_driver_mux_selector);
			track_5_4_chanX_n12 <= track_5_4_chanX_n12_driver_mux_fanins(track_5_4_chanX_n12_driver_mux_selector);
			track_5_4_chanX_n13 <= track_5_4_chanX_n13_driver_mux_fanins(track_5_4_chanX_n13_driver_mux_selector);
			track_5_4_chanX_n14 <= track_5_4_chanX_n14_driver_mux_fanins(track_5_4_chanX_n14_driver_mux_selector);
			track_5_4_chanX_n15 <= track_5_4_chanX_n15_driver_mux_fanins(track_5_4_chanX_n15_driver_mux_selector);
			track_5_4_chanX_n2  <= track_5_4_chanX_n2_driver_mux_fanins(track_5_4_chanX_n2_driver_mux_selector);
			track_5_4_chanX_n3  <= track_5_4_chanX_n3_driver_mux_fanins(track_5_4_chanX_n3_driver_mux_selector);
			track_5_4_chanX_n4  <= track_5_4_chanX_n4_driver_mux_fanins(track_5_4_chanX_n4_driver_mux_selector);
			track_5_4_chanX_n5  <= track_5_4_chanX_n5_driver_mux_fanins(track_5_4_chanX_n5_driver_mux_selector);
			track_5_4_chanX_n6  <= track_5_4_chanX_n6_driver_mux_fanins(track_5_4_chanX_n6_driver_mux_selector);
			track_5_4_chanX_n7  <= track_5_4_chanX_n7_driver_mux_fanins(track_5_4_chanX_n7_driver_mux_selector);
			track_5_4_chanX_n8  <= track_5_4_chanX_n8_driver_mux_fanins(track_5_4_chanX_n8_driver_mux_selector);
			track_5_4_chanX_n9  <= track_5_4_chanX_n9_driver_mux_fanins(track_5_4_chanX_n9_driver_mux_selector);
			track_5_4_chanY_n0  <= track_5_4_chanY_n0_driver_mux_fanins(track_5_4_chanY_n0_driver_mux_selector);
			track_5_4_chanY_n1  <= track_5_4_chanY_n1_driver_mux_fanins(track_5_4_chanY_n1_driver_mux_selector);
			track_5_4_chanY_n10 <= track_5_4_chanY_n10_driver_mux_fanins(track_5_4_chanY_n10_driver_mux_selector);
			track_5_4_chanY_n11 <= track_5_4_chanY_n11_driver_mux_fanins(track_5_4_chanY_n11_driver_mux_selector);
			track_5_4_chanY_n12 <= track_5_4_chanY_n12_driver_mux_fanins(track_5_4_chanY_n12_driver_mux_selector);
			track_5_4_chanY_n13 <= track_5_4_chanY_n13_driver_mux_fanins(track_5_4_chanY_n13_driver_mux_selector);
			track_5_4_chanY_n14 <= track_5_4_chanY_n14_driver_mux_fanins(track_5_4_chanY_n14_driver_mux_selector);
			track_5_4_chanY_n15 <= track_5_4_chanY_n15_driver_mux_fanins(track_5_4_chanY_n15_driver_mux_selector);
			track_5_4_chanY_n2  <= track_5_4_chanY_n2_driver_mux_fanins(track_5_4_chanY_n2_driver_mux_selector);
			track_5_4_chanY_n3  <= track_5_4_chanY_n3_driver_mux_fanins(track_5_4_chanY_n3_driver_mux_selector);
			track_5_4_chanY_n4  <= track_5_4_chanY_n4_driver_mux_fanins(track_5_4_chanY_n4_driver_mux_selector);
			track_5_4_chanY_n5  <= track_5_4_chanY_n5_driver_mux_fanins(track_5_4_chanY_n5_driver_mux_selector);
			track_5_4_chanY_n6  <= track_5_4_chanY_n6_driver_mux_fanins(track_5_4_chanY_n6_driver_mux_selector);
			track_5_4_chanY_n7  <= track_5_4_chanY_n7_driver_mux_fanins(track_5_4_chanY_n7_driver_mux_selector);
			track_5_4_chanY_n8  <= track_5_4_chanY_n8_driver_mux_fanins(track_5_4_chanY_n8_driver_mux_selector);
			track_5_4_chanY_n9  <= track_5_4_chanY_n9_driver_mux_fanins(track_5_4_chanY_n9_driver_mux_selector);
			track_5_5_chanX_n0  <= track_5_5_chanX_n0_driver_mux_fanins(track_5_5_chanX_n0_driver_mux_selector);
			track_5_5_chanX_n1  <= track_5_5_chanX_n1_driver_mux_fanins(track_5_5_chanX_n1_driver_mux_selector);
			track_5_5_chanX_n10 <= track_5_5_chanX_n10_driver_mux_fanins(track_5_5_chanX_n10_driver_mux_selector);
			track_5_5_chanX_n11 <= track_5_5_chanX_n11_driver_mux_fanins(track_5_5_chanX_n11_driver_mux_selector);
			track_5_5_chanX_n12 <= track_5_5_chanX_n12_driver_mux_fanins(track_5_5_chanX_n12_driver_mux_selector);
			track_5_5_chanX_n13 <= track_5_5_chanX_n13_driver_mux_fanins(track_5_5_chanX_n13_driver_mux_selector);
			track_5_5_chanX_n14 <= track_5_5_chanX_n14_driver_mux_fanins(track_5_5_chanX_n14_driver_mux_selector);
			track_5_5_chanX_n15 <= track_5_5_chanX_n15_driver_mux_fanins(track_5_5_chanX_n15_driver_mux_selector);
			track_5_5_chanX_n2  <= track_5_5_chanX_n2_driver_mux_fanins(track_5_5_chanX_n2_driver_mux_selector);
			track_5_5_chanX_n3  <= track_5_5_chanX_n3_driver_mux_fanins(track_5_5_chanX_n3_driver_mux_selector);
			track_5_5_chanX_n4  <= track_5_5_chanX_n4_driver_mux_fanins(track_5_5_chanX_n4_driver_mux_selector);
			track_5_5_chanX_n5  <= track_5_5_chanX_n5_driver_mux_fanins(track_5_5_chanX_n5_driver_mux_selector);
			track_5_5_chanX_n6  <= track_5_5_chanX_n6_driver_mux_fanins(track_5_5_chanX_n6_driver_mux_selector);
			track_5_5_chanX_n7  <= track_5_5_chanX_n7_driver_mux_fanins(track_5_5_chanX_n7_driver_mux_selector);
			track_5_5_chanX_n8  <= track_5_5_chanX_n8_driver_mux_fanins(track_5_5_chanX_n8_driver_mux_selector);
			track_5_5_chanX_n9  <= track_5_5_chanX_n9_driver_mux_fanins(track_5_5_chanX_n9_driver_mux_selector);
			track_5_5_chanY_n0  <= track_5_5_chanY_n0_driver_mux_fanins(track_5_5_chanY_n0_driver_mux_selector);
			track_5_5_chanY_n1  <= track_5_5_chanY_n1_driver_mux_fanins(track_5_5_chanY_n1_driver_mux_selector);
			track_5_5_chanY_n10 <= track_5_5_chanY_n10_driver_mux_fanins(track_5_5_chanY_n10_driver_mux_selector);
			track_5_5_chanY_n11 <= track_5_5_chanY_n11_driver_mux_fanins(track_5_5_chanY_n11_driver_mux_selector);
			track_5_5_chanY_n12 <= track_5_5_chanY_n12_driver_mux_fanins(track_5_5_chanY_n12_driver_mux_selector);
			track_5_5_chanY_n13 <= track_5_5_chanY_n13_driver_mux_fanins(track_5_5_chanY_n13_driver_mux_selector);
			track_5_5_chanY_n14 <= track_5_5_chanY_n14_driver_mux_fanins(track_5_5_chanY_n14_driver_mux_selector);
			track_5_5_chanY_n15 <= track_5_5_chanY_n15_driver_mux_fanins(track_5_5_chanY_n15_driver_mux_selector);
			track_5_5_chanY_n2  <= track_5_5_chanY_n2_driver_mux_fanins(track_5_5_chanY_n2_driver_mux_selector);
			track_5_5_chanY_n3  <= track_5_5_chanY_n3_driver_mux_fanins(track_5_5_chanY_n3_driver_mux_selector);
			track_5_5_chanY_n4  <= track_5_5_chanY_n4_driver_mux_fanins(track_5_5_chanY_n4_driver_mux_selector);
			track_5_5_chanY_n5  <= track_5_5_chanY_n5_driver_mux_fanins(track_5_5_chanY_n5_driver_mux_selector);
			track_5_5_chanY_n6  <= track_5_5_chanY_n6_driver_mux_fanins(track_5_5_chanY_n6_driver_mux_selector);
			track_5_5_chanY_n7  <= track_5_5_chanY_n7_driver_mux_fanins(track_5_5_chanY_n7_driver_mux_selector);
			track_5_5_chanY_n8  <= track_5_5_chanY_n8_driver_mux_fanins(track_5_5_chanY_n8_driver_mux_selector);
			track_5_5_chanY_n9  <= track_5_5_chanY_n9_driver_mux_fanins(track_5_5_chanY_n9_driver_mux_selector);
			track_5_6_chanX_n0  <= track_5_6_chanX_n0_driver_mux_fanins(track_5_6_chanX_n0_driver_mux_selector);
			track_5_6_chanX_n1  <= track_5_6_chanX_n1_driver_mux_fanins(track_5_6_chanX_n1_driver_mux_selector);
			track_5_6_chanX_n10 <= track_5_6_chanX_n10_driver_mux_fanins(track_5_6_chanX_n10_driver_mux_selector);
			track_5_6_chanX_n11 <= track_5_6_chanX_n11_driver_mux_fanins(track_5_6_chanX_n11_driver_mux_selector);
			track_5_6_chanX_n12 <= track_5_6_chanX_n12_driver_mux_fanins(track_5_6_chanX_n12_driver_mux_selector);
			track_5_6_chanX_n13 <= track_5_6_chanX_n13_driver_mux_fanins(track_5_6_chanX_n13_driver_mux_selector);
			track_5_6_chanX_n14 <= track_5_6_chanX_n14_driver_mux_fanins(track_5_6_chanX_n14_driver_mux_selector);
			track_5_6_chanX_n15 <= track_5_6_chanX_n15_driver_mux_fanins(track_5_6_chanX_n15_driver_mux_selector);
			track_5_6_chanX_n2  <= track_5_6_chanX_n2_driver_mux_fanins(track_5_6_chanX_n2_driver_mux_selector);
			track_5_6_chanX_n3  <= track_5_6_chanX_n3_driver_mux_fanins(track_5_6_chanX_n3_driver_mux_selector);
			track_5_6_chanX_n4  <= track_5_6_chanX_n4_driver_mux_fanins(track_5_6_chanX_n4_driver_mux_selector);
			track_5_6_chanX_n5  <= track_5_6_chanX_n5_driver_mux_fanins(track_5_6_chanX_n5_driver_mux_selector);
			track_5_6_chanX_n6  <= track_5_6_chanX_n6_driver_mux_fanins(track_5_6_chanX_n6_driver_mux_selector);
			track_5_6_chanX_n7  <= track_5_6_chanX_n7_driver_mux_fanins(track_5_6_chanX_n7_driver_mux_selector);
			track_5_6_chanX_n8  <= track_5_6_chanX_n8_driver_mux_fanins(track_5_6_chanX_n8_driver_mux_selector);
			track_5_6_chanX_n9  <= track_5_6_chanX_n9_driver_mux_fanins(track_5_6_chanX_n9_driver_mux_selector);
			track_5_6_chanY_n0  <= track_5_6_chanY_n0_driver_mux_fanins(track_5_6_chanY_n0_driver_mux_selector);
			track_5_6_chanY_n1  <= track_5_6_chanY_n1_driver_mux_fanins(track_5_6_chanY_n1_driver_mux_selector);
			track_5_6_chanY_n10 <= track_5_6_chanY_n10_driver_mux_fanins(track_5_6_chanY_n10_driver_mux_selector);
			track_5_6_chanY_n11 <= track_5_6_chanY_n11_driver_mux_fanins(track_5_6_chanY_n11_driver_mux_selector);
			track_5_6_chanY_n12 <= track_5_6_chanY_n12_driver_mux_fanins(track_5_6_chanY_n12_driver_mux_selector);
			track_5_6_chanY_n13 <= track_5_6_chanY_n13_driver_mux_fanins(track_5_6_chanY_n13_driver_mux_selector);
			track_5_6_chanY_n14 <= track_5_6_chanY_n14_driver_mux_fanins(track_5_6_chanY_n14_driver_mux_selector);
			track_5_6_chanY_n15 <= track_5_6_chanY_n15_driver_mux_fanins(track_5_6_chanY_n15_driver_mux_selector);
			track_5_6_chanY_n2  <= track_5_6_chanY_n2_driver_mux_fanins(track_5_6_chanY_n2_driver_mux_selector);
			track_5_6_chanY_n3  <= track_5_6_chanY_n3_driver_mux_fanins(track_5_6_chanY_n3_driver_mux_selector);
			track_5_6_chanY_n4  <= track_5_6_chanY_n4_driver_mux_fanins(track_5_6_chanY_n4_driver_mux_selector);
			track_5_6_chanY_n5  <= track_5_6_chanY_n5_driver_mux_fanins(track_5_6_chanY_n5_driver_mux_selector);
			track_5_6_chanY_n6  <= track_5_6_chanY_n6_driver_mux_fanins(track_5_6_chanY_n6_driver_mux_selector);
			track_5_6_chanY_n7  <= track_5_6_chanY_n7_driver_mux_fanins(track_5_6_chanY_n7_driver_mux_selector);
			track_5_6_chanY_n8  <= track_5_6_chanY_n8_driver_mux_fanins(track_5_6_chanY_n8_driver_mux_selector);
			track_5_6_chanY_n9  <= track_5_6_chanY_n9_driver_mux_fanins(track_5_6_chanY_n9_driver_mux_selector);
			track_6_0_chanX_n0  <= track_6_0_chanX_n0_driver_mux_fanins(track_6_0_chanX_n0_driver_mux_selector);
			track_6_0_chanX_n1  <= track_6_0_chanX_n1_driver_mux_fanins(track_6_0_chanX_n1_driver_mux_selector);
			track_6_0_chanX_n10 <= track_6_0_chanX_n10_driver_mux_fanins(track_6_0_chanX_n10_driver_mux_selector);
			track_6_0_chanX_n11 <= track_6_0_chanX_n11_driver_mux_fanins(track_6_0_chanX_n11_driver_mux_selector);
			track_6_0_chanX_n12 <= track_6_0_chanX_n12_driver_mux_fanins(track_6_0_chanX_n12_driver_mux_selector);
			track_6_0_chanX_n13 <= track_6_0_chanX_n13_driver_mux_fanins(track_6_0_chanX_n13_driver_mux_selector);
			track_6_0_chanX_n14 <= track_6_0_chanX_n14_driver_mux_fanins(track_6_0_chanX_n14_driver_mux_selector);
			track_6_0_chanX_n15 <= track_6_0_chanX_n15_driver_mux_fanins(track_6_0_chanX_n15_driver_mux_selector);
			track_6_0_chanX_n2  <= track_6_0_chanX_n2_driver_mux_fanins(track_6_0_chanX_n2_driver_mux_selector);
			track_6_0_chanX_n3  <= track_6_0_chanX_n3_driver_mux_fanins(track_6_0_chanX_n3_driver_mux_selector);
			track_6_0_chanX_n4  <= track_6_0_chanX_n4_driver_mux_fanins(track_6_0_chanX_n4_driver_mux_selector);
			track_6_0_chanX_n5  <= track_6_0_chanX_n5_driver_mux_fanins(track_6_0_chanX_n5_driver_mux_selector);
			track_6_0_chanX_n6  <= track_6_0_chanX_n6_driver_mux_fanins(track_6_0_chanX_n6_driver_mux_selector);
			track_6_0_chanX_n7  <= track_6_0_chanX_n7_driver_mux_fanins(track_6_0_chanX_n7_driver_mux_selector);
			track_6_0_chanX_n8  <= track_6_0_chanX_n8_driver_mux_fanins(track_6_0_chanX_n8_driver_mux_selector);
			track_6_0_chanX_n9  <= track_6_0_chanX_n9_driver_mux_fanins(track_6_0_chanX_n9_driver_mux_selector);
			track_6_1_chanX_n0  <= track_6_1_chanX_n0_driver_mux_fanins(track_6_1_chanX_n0_driver_mux_selector);
			track_6_1_chanX_n1  <= track_6_1_chanX_n1_driver_mux_fanins(track_6_1_chanX_n1_driver_mux_selector);
			track_6_1_chanX_n10 <= track_6_1_chanX_n10_driver_mux_fanins(track_6_1_chanX_n10_driver_mux_selector);
			track_6_1_chanX_n11 <= track_6_1_chanX_n11_driver_mux_fanins(track_6_1_chanX_n11_driver_mux_selector);
			track_6_1_chanX_n12 <= track_6_1_chanX_n12_driver_mux_fanins(track_6_1_chanX_n12_driver_mux_selector);
			track_6_1_chanX_n13 <= track_6_1_chanX_n13_driver_mux_fanins(track_6_1_chanX_n13_driver_mux_selector);
			track_6_1_chanX_n14 <= track_6_1_chanX_n14_driver_mux_fanins(track_6_1_chanX_n14_driver_mux_selector);
			track_6_1_chanX_n15 <= track_6_1_chanX_n15_driver_mux_fanins(track_6_1_chanX_n15_driver_mux_selector);
			track_6_1_chanX_n2  <= track_6_1_chanX_n2_driver_mux_fanins(track_6_1_chanX_n2_driver_mux_selector);
			track_6_1_chanX_n3  <= track_6_1_chanX_n3_driver_mux_fanins(track_6_1_chanX_n3_driver_mux_selector);
			track_6_1_chanX_n4  <= track_6_1_chanX_n4_driver_mux_fanins(track_6_1_chanX_n4_driver_mux_selector);
			track_6_1_chanX_n5  <= track_6_1_chanX_n5_driver_mux_fanins(track_6_1_chanX_n5_driver_mux_selector);
			track_6_1_chanX_n6  <= track_6_1_chanX_n6_driver_mux_fanins(track_6_1_chanX_n6_driver_mux_selector);
			track_6_1_chanX_n7  <= track_6_1_chanX_n7_driver_mux_fanins(track_6_1_chanX_n7_driver_mux_selector);
			track_6_1_chanX_n8  <= track_6_1_chanX_n8_driver_mux_fanins(track_6_1_chanX_n8_driver_mux_selector);
			track_6_1_chanX_n9  <= track_6_1_chanX_n9_driver_mux_fanins(track_6_1_chanX_n9_driver_mux_selector);
			track_6_1_chanY_n0  <= track_6_1_chanY_n0_driver_mux_fanins(track_6_1_chanY_n0_driver_mux_selector);
			track_6_1_chanY_n1  <= track_6_1_chanY_n1_driver_mux_fanins(track_6_1_chanY_n1_driver_mux_selector);
			track_6_1_chanY_n10 <= track_6_1_chanY_n10_driver_mux_fanins(track_6_1_chanY_n10_driver_mux_selector);
			track_6_1_chanY_n11 <= track_6_1_chanY_n11_driver_mux_fanins(track_6_1_chanY_n11_driver_mux_selector);
			track_6_1_chanY_n12 <= track_6_1_chanY_n12_driver_mux_fanins(track_6_1_chanY_n12_driver_mux_selector);
			track_6_1_chanY_n13 <= track_6_1_chanY_n13_driver_mux_fanins(track_6_1_chanY_n13_driver_mux_selector);
			track_6_1_chanY_n14 <= track_6_1_chanY_n14_driver_mux_fanins(track_6_1_chanY_n14_driver_mux_selector);
			track_6_1_chanY_n15 <= track_6_1_chanY_n15_driver_mux_fanins(track_6_1_chanY_n15_driver_mux_selector);
			track_6_1_chanY_n2  <= track_6_1_chanY_n2_driver_mux_fanins(track_6_1_chanY_n2_driver_mux_selector);
			track_6_1_chanY_n3  <= track_6_1_chanY_n3_driver_mux_fanins(track_6_1_chanY_n3_driver_mux_selector);
			track_6_1_chanY_n4  <= track_6_1_chanY_n4_driver_mux_fanins(track_6_1_chanY_n4_driver_mux_selector);
			track_6_1_chanY_n5  <= track_6_1_chanY_n5_driver_mux_fanins(track_6_1_chanY_n5_driver_mux_selector);
			track_6_1_chanY_n6  <= track_6_1_chanY_n6_driver_mux_fanins(track_6_1_chanY_n6_driver_mux_selector);
			track_6_1_chanY_n7  <= track_6_1_chanY_n7_driver_mux_fanins(track_6_1_chanY_n7_driver_mux_selector);
			track_6_1_chanY_n8  <= track_6_1_chanY_n8_driver_mux_fanins(track_6_1_chanY_n8_driver_mux_selector);
			track_6_1_chanY_n9  <= track_6_1_chanY_n9_driver_mux_fanins(track_6_1_chanY_n9_driver_mux_selector);
			track_6_2_chanX_n0  <= track_6_2_chanX_n0_driver_mux_fanins(track_6_2_chanX_n0_driver_mux_selector);
			track_6_2_chanX_n1  <= track_6_2_chanX_n1_driver_mux_fanins(track_6_2_chanX_n1_driver_mux_selector);
			track_6_2_chanX_n10 <= track_6_2_chanX_n10_driver_mux_fanins(track_6_2_chanX_n10_driver_mux_selector);
			track_6_2_chanX_n11 <= track_6_2_chanX_n11_driver_mux_fanins(track_6_2_chanX_n11_driver_mux_selector);
			track_6_2_chanX_n12 <= track_6_2_chanX_n12_driver_mux_fanins(track_6_2_chanX_n12_driver_mux_selector);
			track_6_2_chanX_n13 <= track_6_2_chanX_n13_driver_mux_fanins(track_6_2_chanX_n13_driver_mux_selector);
			track_6_2_chanX_n14 <= track_6_2_chanX_n14_driver_mux_fanins(track_6_2_chanX_n14_driver_mux_selector);
			track_6_2_chanX_n15 <= track_6_2_chanX_n15_driver_mux_fanins(track_6_2_chanX_n15_driver_mux_selector);
			track_6_2_chanX_n2  <= track_6_2_chanX_n2_driver_mux_fanins(track_6_2_chanX_n2_driver_mux_selector);
			track_6_2_chanX_n3  <= track_6_2_chanX_n3_driver_mux_fanins(track_6_2_chanX_n3_driver_mux_selector);
			track_6_2_chanX_n4  <= track_6_2_chanX_n4_driver_mux_fanins(track_6_2_chanX_n4_driver_mux_selector);
			track_6_2_chanX_n5  <= track_6_2_chanX_n5_driver_mux_fanins(track_6_2_chanX_n5_driver_mux_selector);
			track_6_2_chanX_n6  <= track_6_2_chanX_n6_driver_mux_fanins(track_6_2_chanX_n6_driver_mux_selector);
			track_6_2_chanX_n7  <= track_6_2_chanX_n7_driver_mux_fanins(track_6_2_chanX_n7_driver_mux_selector);
			track_6_2_chanX_n8  <= track_6_2_chanX_n8_driver_mux_fanins(track_6_2_chanX_n8_driver_mux_selector);
			track_6_2_chanX_n9  <= track_6_2_chanX_n9_driver_mux_fanins(track_6_2_chanX_n9_driver_mux_selector);
			track_6_2_chanY_n0  <= track_6_2_chanY_n0_driver_mux_fanins(track_6_2_chanY_n0_driver_mux_selector);
			track_6_2_chanY_n1  <= track_6_2_chanY_n1_driver_mux_fanins(track_6_2_chanY_n1_driver_mux_selector);
			track_6_2_chanY_n10 <= track_6_2_chanY_n10_driver_mux_fanins(track_6_2_chanY_n10_driver_mux_selector);
			track_6_2_chanY_n11 <= track_6_2_chanY_n11_driver_mux_fanins(track_6_2_chanY_n11_driver_mux_selector);
			track_6_2_chanY_n12 <= track_6_2_chanY_n12_driver_mux_fanins(track_6_2_chanY_n12_driver_mux_selector);
			track_6_2_chanY_n13 <= track_6_2_chanY_n13_driver_mux_fanins(track_6_2_chanY_n13_driver_mux_selector);
			track_6_2_chanY_n14 <= track_6_2_chanY_n14_driver_mux_fanins(track_6_2_chanY_n14_driver_mux_selector);
			track_6_2_chanY_n15 <= track_6_2_chanY_n15_driver_mux_fanins(track_6_2_chanY_n15_driver_mux_selector);
			track_6_2_chanY_n2  <= track_6_2_chanY_n2_driver_mux_fanins(track_6_2_chanY_n2_driver_mux_selector);
			track_6_2_chanY_n3  <= track_6_2_chanY_n3_driver_mux_fanins(track_6_2_chanY_n3_driver_mux_selector);
			track_6_2_chanY_n4  <= track_6_2_chanY_n4_driver_mux_fanins(track_6_2_chanY_n4_driver_mux_selector);
			track_6_2_chanY_n5  <= track_6_2_chanY_n5_driver_mux_fanins(track_6_2_chanY_n5_driver_mux_selector);
			track_6_2_chanY_n6  <= track_6_2_chanY_n6_driver_mux_fanins(track_6_2_chanY_n6_driver_mux_selector);
			track_6_2_chanY_n7  <= track_6_2_chanY_n7_driver_mux_fanins(track_6_2_chanY_n7_driver_mux_selector);
			track_6_2_chanY_n8  <= track_6_2_chanY_n8_driver_mux_fanins(track_6_2_chanY_n8_driver_mux_selector);
			track_6_2_chanY_n9  <= track_6_2_chanY_n9_driver_mux_fanins(track_6_2_chanY_n9_driver_mux_selector);
			track_6_3_chanX_n0  <= track_6_3_chanX_n0_driver_mux_fanins(track_6_3_chanX_n0_driver_mux_selector);
			track_6_3_chanX_n1  <= track_6_3_chanX_n1_driver_mux_fanins(track_6_3_chanX_n1_driver_mux_selector);
			track_6_3_chanX_n10 <= track_6_3_chanX_n10_driver_mux_fanins(track_6_3_chanX_n10_driver_mux_selector);
			track_6_3_chanX_n11 <= track_6_3_chanX_n11_driver_mux_fanins(track_6_3_chanX_n11_driver_mux_selector);
			track_6_3_chanX_n12 <= track_6_3_chanX_n12_driver_mux_fanins(track_6_3_chanX_n12_driver_mux_selector);
			track_6_3_chanX_n13 <= track_6_3_chanX_n13_driver_mux_fanins(track_6_3_chanX_n13_driver_mux_selector);
			track_6_3_chanX_n14 <= track_6_3_chanX_n14_driver_mux_fanins(track_6_3_chanX_n14_driver_mux_selector);
			track_6_3_chanX_n15 <= track_6_3_chanX_n15_driver_mux_fanins(track_6_3_chanX_n15_driver_mux_selector);
			track_6_3_chanX_n2  <= track_6_3_chanX_n2_driver_mux_fanins(track_6_3_chanX_n2_driver_mux_selector);
			track_6_3_chanX_n3  <= track_6_3_chanX_n3_driver_mux_fanins(track_6_3_chanX_n3_driver_mux_selector);
			track_6_3_chanX_n4  <= track_6_3_chanX_n4_driver_mux_fanins(track_6_3_chanX_n4_driver_mux_selector);
			track_6_3_chanX_n5  <= track_6_3_chanX_n5_driver_mux_fanins(track_6_3_chanX_n5_driver_mux_selector);
			track_6_3_chanX_n6  <= track_6_3_chanX_n6_driver_mux_fanins(track_6_3_chanX_n6_driver_mux_selector);
			track_6_3_chanX_n7  <= track_6_3_chanX_n7_driver_mux_fanins(track_6_3_chanX_n7_driver_mux_selector);
			track_6_3_chanX_n8  <= track_6_3_chanX_n8_driver_mux_fanins(track_6_3_chanX_n8_driver_mux_selector);
			track_6_3_chanX_n9  <= track_6_3_chanX_n9_driver_mux_fanins(track_6_3_chanX_n9_driver_mux_selector);
			track_6_3_chanY_n0  <= track_6_3_chanY_n0_driver_mux_fanins(track_6_3_chanY_n0_driver_mux_selector);
			track_6_3_chanY_n1  <= track_6_3_chanY_n1_driver_mux_fanins(track_6_3_chanY_n1_driver_mux_selector);
			track_6_3_chanY_n10 <= track_6_3_chanY_n10_driver_mux_fanins(track_6_3_chanY_n10_driver_mux_selector);
			track_6_3_chanY_n11 <= track_6_3_chanY_n11_driver_mux_fanins(track_6_3_chanY_n11_driver_mux_selector);
			track_6_3_chanY_n12 <= track_6_3_chanY_n12_driver_mux_fanins(track_6_3_chanY_n12_driver_mux_selector);
			track_6_3_chanY_n13 <= track_6_3_chanY_n13_driver_mux_fanins(track_6_3_chanY_n13_driver_mux_selector);
			track_6_3_chanY_n14 <= track_6_3_chanY_n14_driver_mux_fanins(track_6_3_chanY_n14_driver_mux_selector);
			track_6_3_chanY_n15 <= track_6_3_chanY_n15_driver_mux_fanins(track_6_3_chanY_n15_driver_mux_selector);
			track_6_3_chanY_n2  <= track_6_3_chanY_n2_driver_mux_fanins(track_6_3_chanY_n2_driver_mux_selector);
			track_6_3_chanY_n3  <= track_6_3_chanY_n3_driver_mux_fanins(track_6_3_chanY_n3_driver_mux_selector);
			track_6_3_chanY_n4  <= track_6_3_chanY_n4_driver_mux_fanins(track_6_3_chanY_n4_driver_mux_selector);
			track_6_3_chanY_n5  <= track_6_3_chanY_n5_driver_mux_fanins(track_6_3_chanY_n5_driver_mux_selector);
			track_6_3_chanY_n6  <= track_6_3_chanY_n6_driver_mux_fanins(track_6_3_chanY_n6_driver_mux_selector);
			track_6_3_chanY_n7  <= track_6_3_chanY_n7_driver_mux_fanins(track_6_3_chanY_n7_driver_mux_selector);
			track_6_3_chanY_n8  <= track_6_3_chanY_n8_driver_mux_fanins(track_6_3_chanY_n8_driver_mux_selector);
			track_6_3_chanY_n9  <= track_6_3_chanY_n9_driver_mux_fanins(track_6_3_chanY_n9_driver_mux_selector);
			track_6_4_chanX_n0  <= track_6_4_chanX_n0_driver_mux_fanins(track_6_4_chanX_n0_driver_mux_selector);
			track_6_4_chanX_n1  <= track_6_4_chanX_n1_driver_mux_fanins(track_6_4_chanX_n1_driver_mux_selector);
			track_6_4_chanX_n10 <= track_6_4_chanX_n10_driver_mux_fanins(track_6_4_chanX_n10_driver_mux_selector);
			track_6_4_chanX_n11 <= track_6_4_chanX_n11_driver_mux_fanins(track_6_4_chanX_n11_driver_mux_selector);
			track_6_4_chanX_n12 <= track_6_4_chanX_n12_driver_mux_fanins(track_6_4_chanX_n12_driver_mux_selector);
			track_6_4_chanX_n13 <= track_6_4_chanX_n13_driver_mux_fanins(track_6_4_chanX_n13_driver_mux_selector);
			track_6_4_chanX_n14 <= track_6_4_chanX_n14_driver_mux_fanins(track_6_4_chanX_n14_driver_mux_selector);
			track_6_4_chanX_n15 <= track_6_4_chanX_n15_driver_mux_fanins(track_6_4_chanX_n15_driver_mux_selector);
			track_6_4_chanX_n2  <= track_6_4_chanX_n2_driver_mux_fanins(track_6_4_chanX_n2_driver_mux_selector);
			track_6_4_chanX_n3  <= track_6_4_chanX_n3_driver_mux_fanins(track_6_4_chanX_n3_driver_mux_selector);
			track_6_4_chanX_n4  <= track_6_4_chanX_n4_driver_mux_fanins(track_6_4_chanX_n4_driver_mux_selector);
			track_6_4_chanX_n5  <= track_6_4_chanX_n5_driver_mux_fanins(track_6_4_chanX_n5_driver_mux_selector);
			track_6_4_chanX_n6  <= track_6_4_chanX_n6_driver_mux_fanins(track_6_4_chanX_n6_driver_mux_selector);
			track_6_4_chanX_n7  <= track_6_4_chanX_n7_driver_mux_fanins(track_6_4_chanX_n7_driver_mux_selector);
			track_6_4_chanX_n8  <= track_6_4_chanX_n8_driver_mux_fanins(track_6_4_chanX_n8_driver_mux_selector);
			track_6_4_chanX_n9  <= track_6_4_chanX_n9_driver_mux_fanins(track_6_4_chanX_n9_driver_mux_selector);
			track_6_4_chanY_n0  <= track_6_4_chanY_n0_driver_mux_fanins(track_6_4_chanY_n0_driver_mux_selector);
			track_6_4_chanY_n1  <= track_6_4_chanY_n1_driver_mux_fanins(track_6_4_chanY_n1_driver_mux_selector);
			track_6_4_chanY_n10 <= track_6_4_chanY_n10_driver_mux_fanins(track_6_4_chanY_n10_driver_mux_selector);
			track_6_4_chanY_n11 <= track_6_4_chanY_n11_driver_mux_fanins(track_6_4_chanY_n11_driver_mux_selector);
			track_6_4_chanY_n12 <= track_6_4_chanY_n12_driver_mux_fanins(track_6_4_chanY_n12_driver_mux_selector);
			track_6_4_chanY_n13 <= track_6_4_chanY_n13_driver_mux_fanins(track_6_4_chanY_n13_driver_mux_selector);
			track_6_4_chanY_n14 <= track_6_4_chanY_n14_driver_mux_fanins(track_6_4_chanY_n14_driver_mux_selector);
			track_6_4_chanY_n15 <= track_6_4_chanY_n15_driver_mux_fanins(track_6_4_chanY_n15_driver_mux_selector);
			track_6_4_chanY_n2  <= track_6_4_chanY_n2_driver_mux_fanins(track_6_4_chanY_n2_driver_mux_selector);
			track_6_4_chanY_n3  <= track_6_4_chanY_n3_driver_mux_fanins(track_6_4_chanY_n3_driver_mux_selector);
			track_6_4_chanY_n4  <= track_6_4_chanY_n4_driver_mux_fanins(track_6_4_chanY_n4_driver_mux_selector);
			track_6_4_chanY_n5  <= track_6_4_chanY_n5_driver_mux_fanins(track_6_4_chanY_n5_driver_mux_selector);
			track_6_4_chanY_n6  <= track_6_4_chanY_n6_driver_mux_fanins(track_6_4_chanY_n6_driver_mux_selector);
			track_6_4_chanY_n7  <= track_6_4_chanY_n7_driver_mux_fanins(track_6_4_chanY_n7_driver_mux_selector);
			track_6_4_chanY_n8  <= track_6_4_chanY_n8_driver_mux_fanins(track_6_4_chanY_n8_driver_mux_selector);
			track_6_4_chanY_n9  <= track_6_4_chanY_n9_driver_mux_fanins(track_6_4_chanY_n9_driver_mux_selector);
			track_6_5_chanX_n0  <= track_6_5_chanX_n0_driver_mux_fanins(track_6_5_chanX_n0_driver_mux_selector);
			track_6_5_chanX_n1  <= track_6_5_chanX_n1_driver_mux_fanins(track_6_5_chanX_n1_driver_mux_selector);
			track_6_5_chanX_n10 <= track_6_5_chanX_n10_driver_mux_fanins(track_6_5_chanX_n10_driver_mux_selector);
			track_6_5_chanX_n11 <= track_6_5_chanX_n11_driver_mux_fanins(track_6_5_chanX_n11_driver_mux_selector);
			track_6_5_chanX_n12 <= track_6_5_chanX_n12_driver_mux_fanins(track_6_5_chanX_n12_driver_mux_selector);
			track_6_5_chanX_n13 <= track_6_5_chanX_n13_driver_mux_fanins(track_6_5_chanX_n13_driver_mux_selector);
			track_6_5_chanX_n14 <= track_6_5_chanX_n14_driver_mux_fanins(track_6_5_chanX_n14_driver_mux_selector);
			track_6_5_chanX_n15 <= track_6_5_chanX_n15_driver_mux_fanins(track_6_5_chanX_n15_driver_mux_selector);
			track_6_5_chanX_n2  <= track_6_5_chanX_n2_driver_mux_fanins(track_6_5_chanX_n2_driver_mux_selector);
			track_6_5_chanX_n3  <= track_6_5_chanX_n3_driver_mux_fanins(track_6_5_chanX_n3_driver_mux_selector);
			track_6_5_chanX_n4  <= track_6_5_chanX_n4_driver_mux_fanins(track_6_5_chanX_n4_driver_mux_selector);
			track_6_5_chanX_n5  <= track_6_5_chanX_n5_driver_mux_fanins(track_6_5_chanX_n5_driver_mux_selector);
			track_6_5_chanX_n6  <= track_6_5_chanX_n6_driver_mux_fanins(track_6_5_chanX_n6_driver_mux_selector);
			track_6_5_chanX_n7  <= track_6_5_chanX_n7_driver_mux_fanins(track_6_5_chanX_n7_driver_mux_selector);
			track_6_5_chanX_n8  <= track_6_5_chanX_n8_driver_mux_fanins(track_6_5_chanX_n8_driver_mux_selector);
			track_6_5_chanX_n9  <= track_6_5_chanX_n9_driver_mux_fanins(track_6_5_chanX_n9_driver_mux_selector);
			track_6_5_chanY_n0  <= track_6_5_chanY_n0_driver_mux_fanins(track_6_5_chanY_n0_driver_mux_selector);
			track_6_5_chanY_n1  <= track_6_5_chanY_n1_driver_mux_fanins(track_6_5_chanY_n1_driver_mux_selector);
			track_6_5_chanY_n10 <= track_6_5_chanY_n10_driver_mux_fanins(track_6_5_chanY_n10_driver_mux_selector);
			track_6_5_chanY_n11 <= track_6_5_chanY_n11_driver_mux_fanins(track_6_5_chanY_n11_driver_mux_selector);
			track_6_5_chanY_n12 <= track_6_5_chanY_n12_driver_mux_fanins(track_6_5_chanY_n12_driver_mux_selector);
			track_6_5_chanY_n13 <= track_6_5_chanY_n13_driver_mux_fanins(track_6_5_chanY_n13_driver_mux_selector);
			track_6_5_chanY_n14 <= track_6_5_chanY_n14_driver_mux_fanins(track_6_5_chanY_n14_driver_mux_selector);
			track_6_5_chanY_n15 <= track_6_5_chanY_n15_driver_mux_fanins(track_6_5_chanY_n15_driver_mux_selector);
			track_6_5_chanY_n2  <= track_6_5_chanY_n2_driver_mux_fanins(track_6_5_chanY_n2_driver_mux_selector);
			track_6_5_chanY_n3  <= track_6_5_chanY_n3_driver_mux_fanins(track_6_5_chanY_n3_driver_mux_selector);
			track_6_5_chanY_n4  <= track_6_5_chanY_n4_driver_mux_fanins(track_6_5_chanY_n4_driver_mux_selector);
			track_6_5_chanY_n5  <= track_6_5_chanY_n5_driver_mux_fanins(track_6_5_chanY_n5_driver_mux_selector);
			track_6_5_chanY_n6  <= track_6_5_chanY_n6_driver_mux_fanins(track_6_5_chanY_n6_driver_mux_selector);
			track_6_5_chanY_n7  <= track_6_5_chanY_n7_driver_mux_fanins(track_6_5_chanY_n7_driver_mux_selector);
			track_6_5_chanY_n8  <= track_6_5_chanY_n8_driver_mux_fanins(track_6_5_chanY_n8_driver_mux_selector);
			track_6_5_chanY_n9  <= track_6_5_chanY_n9_driver_mux_fanins(track_6_5_chanY_n9_driver_mux_selector);
			track_6_6_chanX_n0  <= track_6_6_chanX_n0_driver_mux_fanins(track_6_6_chanX_n0_driver_mux_selector);
			track_6_6_chanX_n1  <= track_6_6_chanX_n1_driver_mux_fanins(track_6_6_chanX_n1_driver_mux_selector);
			track_6_6_chanX_n10 <= track_6_6_chanX_n10_driver_mux_fanins(track_6_6_chanX_n10_driver_mux_selector);
			track_6_6_chanX_n11 <= track_6_6_chanX_n11_driver_mux_fanins(track_6_6_chanX_n11_driver_mux_selector);
			track_6_6_chanX_n12 <= track_6_6_chanX_n12_driver_mux_fanins(track_6_6_chanX_n12_driver_mux_selector);
			track_6_6_chanX_n13 <= track_6_6_chanX_n13_driver_mux_fanins(track_6_6_chanX_n13_driver_mux_selector);
			track_6_6_chanX_n14 <= track_6_6_chanX_n14_driver_mux_fanins(track_6_6_chanX_n14_driver_mux_selector);
			track_6_6_chanX_n15 <= track_6_6_chanX_n15_driver_mux_fanins(track_6_6_chanX_n15_driver_mux_selector);
			track_6_6_chanX_n2  <= track_6_6_chanX_n2_driver_mux_fanins(track_6_6_chanX_n2_driver_mux_selector);
			track_6_6_chanX_n3  <= track_6_6_chanX_n3_driver_mux_fanins(track_6_6_chanX_n3_driver_mux_selector);
			track_6_6_chanX_n4  <= track_6_6_chanX_n4_driver_mux_fanins(track_6_6_chanX_n4_driver_mux_selector);
			track_6_6_chanX_n5  <= track_6_6_chanX_n5_driver_mux_fanins(track_6_6_chanX_n5_driver_mux_selector);
			track_6_6_chanX_n6  <= track_6_6_chanX_n6_driver_mux_fanins(track_6_6_chanX_n6_driver_mux_selector);
			track_6_6_chanX_n7  <= track_6_6_chanX_n7_driver_mux_fanins(track_6_6_chanX_n7_driver_mux_selector);
			track_6_6_chanX_n8  <= track_6_6_chanX_n8_driver_mux_fanins(track_6_6_chanX_n8_driver_mux_selector);
			track_6_6_chanX_n9  <= track_6_6_chanX_n9_driver_mux_fanins(track_6_6_chanX_n9_driver_mux_selector);
			track_6_6_chanY_n0  <= track_6_6_chanY_n0_driver_mux_fanins(track_6_6_chanY_n0_driver_mux_selector);
			track_6_6_chanY_n1  <= track_6_6_chanY_n1_driver_mux_fanins(track_6_6_chanY_n1_driver_mux_selector);
			track_6_6_chanY_n10 <= track_6_6_chanY_n10_driver_mux_fanins(track_6_6_chanY_n10_driver_mux_selector);
			track_6_6_chanY_n11 <= track_6_6_chanY_n11_driver_mux_fanins(track_6_6_chanY_n11_driver_mux_selector);
			track_6_6_chanY_n12 <= track_6_6_chanY_n12_driver_mux_fanins(track_6_6_chanY_n12_driver_mux_selector);
			track_6_6_chanY_n13 <= track_6_6_chanY_n13_driver_mux_fanins(track_6_6_chanY_n13_driver_mux_selector);
			track_6_6_chanY_n14 <= track_6_6_chanY_n14_driver_mux_fanins(track_6_6_chanY_n14_driver_mux_selector);
			track_6_6_chanY_n15 <= track_6_6_chanY_n15_driver_mux_fanins(track_6_6_chanY_n15_driver_mux_selector);
			track_6_6_chanY_n2  <= track_6_6_chanY_n2_driver_mux_fanins(track_6_6_chanY_n2_driver_mux_selector);
			track_6_6_chanY_n3  <= track_6_6_chanY_n3_driver_mux_fanins(track_6_6_chanY_n3_driver_mux_selector);
			track_6_6_chanY_n4  <= track_6_6_chanY_n4_driver_mux_fanins(track_6_6_chanY_n4_driver_mux_selector);
			track_6_6_chanY_n5  <= track_6_6_chanY_n5_driver_mux_fanins(track_6_6_chanY_n5_driver_mux_selector);
			track_6_6_chanY_n6  <= track_6_6_chanY_n6_driver_mux_fanins(track_6_6_chanY_n6_driver_mux_selector);
			track_6_6_chanY_n7  <= track_6_6_chanY_n7_driver_mux_fanins(track_6_6_chanY_n7_driver_mux_selector);
			track_6_6_chanY_n8  <= track_6_6_chanY_n8_driver_mux_fanins(track_6_6_chanY_n8_driver_mux_selector);
			track_6_6_chanY_n9  <= track_6_6_chanY_n9_driver_mux_fanins(track_6_6_chanY_n9_driver_mux_selector);
			track_7_0_chanX_n0  <= track_7_0_chanX_n0_driver_mux_fanins(track_7_0_chanX_n0_driver_mux_selector);
			track_7_0_chanX_n1  <= track_7_0_chanX_n1_driver_mux_fanins(track_7_0_chanX_n1_driver_mux_selector);
			track_7_0_chanX_n10 <= track_7_0_chanX_n10_driver_mux_fanins(track_7_0_chanX_n10_driver_mux_selector);
			track_7_0_chanX_n11 <= track_7_0_chanX_n11_driver_mux_fanins(track_7_0_chanX_n11_driver_mux_selector);
			track_7_0_chanX_n12 <= track_7_0_chanX_n12_driver_mux_fanins(track_7_0_chanX_n12_driver_mux_selector);
			track_7_0_chanX_n13 <= track_7_0_chanX_n13_driver_mux_fanins(track_7_0_chanX_n13_driver_mux_selector);
			track_7_0_chanX_n14 <= track_7_0_chanX_n14_driver_mux_fanins(track_7_0_chanX_n14_driver_mux_selector);
			track_7_0_chanX_n15 <= track_7_0_chanX_n15_driver_mux_fanins(track_7_0_chanX_n15_driver_mux_selector);
			track_7_0_chanX_n2  <= track_7_0_chanX_n2_driver_mux_fanins(track_7_0_chanX_n2_driver_mux_selector);
			track_7_0_chanX_n3  <= track_7_0_chanX_n3_driver_mux_fanins(track_7_0_chanX_n3_driver_mux_selector);
			track_7_0_chanX_n4  <= track_7_0_chanX_n4_driver_mux_fanins(track_7_0_chanX_n4_driver_mux_selector);
			track_7_0_chanX_n5  <= track_7_0_chanX_n5_driver_mux_fanins(track_7_0_chanX_n5_driver_mux_selector);
			track_7_0_chanX_n6  <= track_7_0_chanX_n6_driver_mux_fanins(track_7_0_chanX_n6_driver_mux_selector);
			track_7_0_chanX_n7  <= track_7_0_chanX_n7_driver_mux_fanins(track_7_0_chanX_n7_driver_mux_selector);
			track_7_0_chanX_n8  <= track_7_0_chanX_n8_driver_mux_fanins(track_7_0_chanX_n8_driver_mux_selector);
			track_7_0_chanX_n9  <= track_7_0_chanX_n9_driver_mux_fanins(track_7_0_chanX_n9_driver_mux_selector);
			track_7_1_chanX_n0  <= track_7_1_chanX_n0_driver_mux_fanins(track_7_1_chanX_n0_driver_mux_selector);
			track_7_1_chanX_n1  <= track_7_1_chanX_n1_driver_mux_fanins(track_7_1_chanX_n1_driver_mux_selector);
			track_7_1_chanX_n10 <= track_7_1_chanX_n10_driver_mux_fanins(track_7_1_chanX_n10_driver_mux_selector);
			track_7_1_chanX_n11 <= track_7_1_chanX_n11_driver_mux_fanins(track_7_1_chanX_n11_driver_mux_selector);
			track_7_1_chanX_n12 <= track_7_1_chanX_n12_driver_mux_fanins(track_7_1_chanX_n12_driver_mux_selector);
			track_7_1_chanX_n13 <= track_7_1_chanX_n13_driver_mux_fanins(track_7_1_chanX_n13_driver_mux_selector);
			track_7_1_chanX_n14 <= track_7_1_chanX_n14_driver_mux_fanins(track_7_1_chanX_n14_driver_mux_selector);
			track_7_1_chanX_n15 <= track_7_1_chanX_n15_driver_mux_fanins(track_7_1_chanX_n15_driver_mux_selector);
			track_7_1_chanX_n2  <= track_7_1_chanX_n2_driver_mux_fanins(track_7_1_chanX_n2_driver_mux_selector);
			track_7_1_chanX_n3  <= track_7_1_chanX_n3_driver_mux_fanins(track_7_1_chanX_n3_driver_mux_selector);
			track_7_1_chanX_n4  <= track_7_1_chanX_n4_driver_mux_fanins(track_7_1_chanX_n4_driver_mux_selector);
			track_7_1_chanX_n5  <= track_7_1_chanX_n5_driver_mux_fanins(track_7_1_chanX_n5_driver_mux_selector);
			track_7_1_chanX_n6  <= track_7_1_chanX_n6_driver_mux_fanins(track_7_1_chanX_n6_driver_mux_selector);
			track_7_1_chanX_n7  <= track_7_1_chanX_n7_driver_mux_fanins(track_7_1_chanX_n7_driver_mux_selector);
			track_7_1_chanX_n8  <= track_7_1_chanX_n8_driver_mux_fanins(track_7_1_chanX_n8_driver_mux_selector);
			track_7_1_chanX_n9  <= track_7_1_chanX_n9_driver_mux_fanins(track_7_1_chanX_n9_driver_mux_selector);
			track_7_1_chanY_n0  <= track_7_1_chanY_n0_driver_mux_fanins(track_7_1_chanY_n0_driver_mux_selector);
			track_7_1_chanY_n1  <= track_7_1_chanY_n1_driver_mux_fanins(track_7_1_chanY_n1_driver_mux_selector);
			track_7_1_chanY_n10 <= track_7_1_chanY_n10_driver_mux_fanins(track_7_1_chanY_n10_driver_mux_selector);
			track_7_1_chanY_n11 <= track_7_1_chanY_n11_driver_mux_fanins(track_7_1_chanY_n11_driver_mux_selector);
			track_7_1_chanY_n12 <= track_7_1_chanY_n12_driver_mux_fanins(track_7_1_chanY_n12_driver_mux_selector);
			track_7_1_chanY_n13 <= track_7_1_chanY_n13_driver_mux_fanins(track_7_1_chanY_n13_driver_mux_selector);
			track_7_1_chanY_n14 <= track_7_1_chanY_n14_driver_mux_fanins(track_7_1_chanY_n14_driver_mux_selector);
			track_7_1_chanY_n15 <= track_7_1_chanY_n15_driver_mux_fanins(track_7_1_chanY_n15_driver_mux_selector);
			track_7_1_chanY_n2  <= track_7_1_chanY_n2_driver_mux_fanins(track_7_1_chanY_n2_driver_mux_selector);
			track_7_1_chanY_n3  <= track_7_1_chanY_n3_driver_mux_fanins(track_7_1_chanY_n3_driver_mux_selector);
			track_7_1_chanY_n4  <= track_7_1_chanY_n4_driver_mux_fanins(track_7_1_chanY_n4_driver_mux_selector);
			track_7_1_chanY_n5  <= track_7_1_chanY_n5_driver_mux_fanins(track_7_1_chanY_n5_driver_mux_selector);
			track_7_1_chanY_n6  <= track_7_1_chanY_n6_driver_mux_fanins(track_7_1_chanY_n6_driver_mux_selector);
			track_7_1_chanY_n7  <= track_7_1_chanY_n7_driver_mux_fanins(track_7_1_chanY_n7_driver_mux_selector);
			track_7_1_chanY_n8  <= track_7_1_chanY_n8_driver_mux_fanins(track_7_1_chanY_n8_driver_mux_selector);
			track_7_1_chanY_n9  <= track_7_1_chanY_n9_driver_mux_fanins(track_7_1_chanY_n9_driver_mux_selector);
			track_7_2_chanX_n0  <= track_7_2_chanX_n0_driver_mux_fanins(track_7_2_chanX_n0_driver_mux_selector);
			track_7_2_chanX_n1  <= track_7_2_chanX_n1_driver_mux_fanins(track_7_2_chanX_n1_driver_mux_selector);
			track_7_2_chanX_n10 <= track_7_2_chanX_n10_driver_mux_fanins(track_7_2_chanX_n10_driver_mux_selector);
			track_7_2_chanX_n11 <= track_7_2_chanX_n11_driver_mux_fanins(track_7_2_chanX_n11_driver_mux_selector);
			track_7_2_chanX_n12 <= track_7_2_chanX_n12_driver_mux_fanins(track_7_2_chanX_n12_driver_mux_selector);
			track_7_2_chanX_n13 <= track_7_2_chanX_n13_driver_mux_fanins(track_7_2_chanX_n13_driver_mux_selector);
			track_7_2_chanX_n14 <= track_7_2_chanX_n14_driver_mux_fanins(track_7_2_chanX_n14_driver_mux_selector);
			track_7_2_chanX_n15 <= track_7_2_chanX_n15_driver_mux_fanins(track_7_2_chanX_n15_driver_mux_selector);
			track_7_2_chanX_n2  <= track_7_2_chanX_n2_driver_mux_fanins(track_7_2_chanX_n2_driver_mux_selector);
			track_7_2_chanX_n3  <= track_7_2_chanX_n3_driver_mux_fanins(track_7_2_chanX_n3_driver_mux_selector);
			track_7_2_chanX_n4  <= track_7_2_chanX_n4_driver_mux_fanins(track_7_2_chanX_n4_driver_mux_selector);
			track_7_2_chanX_n5  <= track_7_2_chanX_n5_driver_mux_fanins(track_7_2_chanX_n5_driver_mux_selector);
			track_7_2_chanX_n6  <= track_7_2_chanX_n6_driver_mux_fanins(track_7_2_chanX_n6_driver_mux_selector);
			track_7_2_chanX_n7  <= track_7_2_chanX_n7_driver_mux_fanins(track_7_2_chanX_n7_driver_mux_selector);
			track_7_2_chanX_n8  <= track_7_2_chanX_n8_driver_mux_fanins(track_7_2_chanX_n8_driver_mux_selector);
			track_7_2_chanX_n9  <= track_7_2_chanX_n9_driver_mux_fanins(track_7_2_chanX_n9_driver_mux_selector);
			track_7_2_chanY_n0  <= track_7_2_chanY_n0_driver_mux_fanins(track_7_2_chanY_n0_driver_mux_selector);
			track_7_2_chanY_n1  <= track_7_2_chanY_n1_driver_mux_fanins(track_7_2_chanY_n1_driver_mux_selector);
			track_7_2_chanY_n10 <= track_7_2_chanY_n10_driver_mux_fanins(track_7_2_chanY_n10_driver_mux_selector);
			track_7_2_chanY_n11 <= track_7_2_chanY_n11_driver_mux_fanins(track_7_2_chanY_n11_driver_mux_selector);
			track_7_2_chanY_n12 <= track_7_2_chanY_n12_driver_mux_fanins(track_7_2_chanY_n12_driver_mux_selector);
			track_7_2_chanY_n13 <= track_7_2_chanY_n13_driver_mux_fanins(track_7_2_chanY_n13_driver_mux_selector);
			track_7_2_chanY_n14 <= track_7_2_chanY_n14_driver_mux_fanins(track_7_2_chanY_n14_driver_mux_selector);
			track_7_2_chanY_n15 <= track_7_2_chanY_n15_driver_mux_fanins(track_7_2_chanY_n15_driver_mux_selector);
			track_7_2_chanY_n2  <= track_7_2_chanY_n2_driver_mux_fanins(track_7_2_chanY_n2_driver_mux_selector);
			track_7_2_chanY_n3  <= track_7_2_chanY_n3_driver_mux_fanins(track_7_2_chanY_n3_driver_mux_selector);
			track_7_2_chanY_n4  <= track_7_2_chanY_n4_driver_mux_fanins(track_7_2_chanY_n4_driver_mux_selector);
			track_7_2_chanY_n5  <= track_7_2_chanY_n5_driver_mux_fanins(track_7_2_chanY_n5_driver_mux_selector);
			track_7_2_chanY_n6  <= track_7_2_chanY_n6_driver_mux_fanins(track_7_2_chanY_n6_driver_mux_selector);
			track_7_2_chanY_n7  <= track_7_2_chanY_n7_driver_mux_fanins(track_7_2_chanY_n7_driver_mux_selector);
			track_7_2_chanY_n8  <= track_7_2_chanY_n8_driver_mux_fanins(track_7_2_chanY_n8_driver_mux_selector);
			track_7_2_chanY_n9  <= track_7_2_chanY_n9_driver_mux_fanins(track_7_2_chanY_n9_driver_mux_selector);
			track_7_3_chanX_n0  <= track_7_3_chanX_n0_driver_mux_fanins(track_7_3_chanX_n0_driver_mux_selector);
			track_7_3_chanX_n1  <= track_7_3_chanX_n1_driver_mux_fanins(track_7_3_chanX_n1_driver_mux_selector);
			track_7_3_chanX_n10 <= track_7_3_chanX_n10_driver_mux_fanins(track_7_3_chanX_n10_driver_mux_selector);
			track_7_3_chanX_n11 <= track_7_3_chanX_n11_driver_mux_fanins(track_7_3_chanX_n11_driver_mux_selector);
			track_7_3_chanX_n12 <= track_7_3_chanX_n12_driver_mux_fanins(track_7_3_chanX_n12_driver_mux_selector);
			track_7_3_chanX_n13 <= track_7_3_chanX_n13_driver_mux_fanins(track_7_3_chanX_n13_driver_mux_selector);
			track_7_3_chanX_n14 <= track_7_3_chanX_n14_driver_mux_fanins(track_7_3_chanX_n14_driver_mux_selector);
			track_7_3_chanX_n15 <= track_7_3_chanX_n15_driver_mux_fanins(track_7_3_chanX_n15_driver_mux_selector);
			track_7_3_chanX_n2  <= track_7_3_chanX_n2_driver_mux_fanins(track_7_3_chanX_n2_driver_mux_selector);
			track_7_3_chanX_n3  <= track_7_3_chanX_n3_driver_mux_fanins(track_7_3_chanX_n3_driver_mux_selector);
			track_7_3_chanX_n4  <= track_7_3_chanX_n4_driver_mux_fanins(track_7_3_chanX_n4_driver_mux_selector);
			track_7_3_chanX_n5  <= track_7_3_chanX_n5_driver_mux_fanins(track_7_3_chanX_n5_driver_mux_selector);
			track_7_3_chanX_n6  <= track_7_3_chanX_n6_driver_mux_fanins(track_7_3_chanX_n6_driver_mux_selector);
			track_7_3_chanX_n7  <= track_7_3_chanX_n7_driver_mux_fanins(track_7_3_chanX_n7_driver_mux_selector);
			track_7_3_chanX_n8  <= track_7_3_chanX_n8_driver_mux_fanins(track_7_3_chanX_n8_driver_mux_selector);
			track_7_3_chanX_n9  <= track_7_3_chanX_n9_driver_mux_fanins(track_7_3_chanX_n9_driver_mux_selector);
			track_7_3_chanY_n0  <= track_7_3_chanY_n0_driver_mux_fanins(track_7_3_chanY_n0_driver_mux_selector);
			track_7_3_chanY_n1  <= track_7_3_chanY_n1_driver_mux_fanins(track_7_3_chanY_n1_driver_mux_selector);
			track_7_3_chanY_n10 <= track_7_3_chanY_n10_driver_mux_fanins(track_7_3_chanY_n10_driver_mux_selector);
			track_7_3_chanY_n11 <= track_7_3_chanY_n11_driver_mux_fanins(track_7_3_chanY_n11_driver_mux_selector);
			track_7_3_chanY_n12 <= track_7_3_chanY_n12_driver_mux_fanins(track_7_3_chanY_n12_driver_mux_selector);
			track_7_3_chanY_n13 <= track_7_3_chanY_n13_driver_mux_fanins(track_7_3_chanY_n13_driver_mux_selector);
			track_7_3_chanY_n14 <= track_7_3_chanY_n14_driver_mux_fanins(track_7_3_chanY_n14_driver_mux_selector);
			track_7_3_chanY_n15 <= track_7_3_chanY_n15_driver_mux_fanins(track_7_3_chanY_n15_driver_mux_selector);
			track_7_3_chanY_n2  <= track_7_3_chanY_n2_driver_mux_fanins(track_7_3_chanY_n2_driver_mux_selector);
			track_7_3_chanY_n3  <= track_7_3_chanY_n3_driver_mux_fanins(track_7_3_chanY_n3_driver_mux_selector);
			track_7_3_chanY_n4  <= track_7_3_chanY_n4_driver_mux_fanins(track_7_3_chanY_n4_driver_mux_selector);
			track_7_3_chanY_n5  <= track_7_3_chanY_n5_driver_mux_fanins(track_7_3_chanY_n5_driver_mux_selector);
			track_7_3_chanY_n6  <= track_7_3_chanY_n6_driver_mux_fanins(track_7_3_chanY_n6_driver_mux_selector);
			track_7_3_chanY_n7  <= track_7_3_chanY_n7_driver_mux_fanins(track_7_3_chanY_n7_driver_mux_selector);
			track_7_3_chanY_n8  <= track_7_3_chanY_n8_driver_mux_fanins(track_7_3_chanY_n8_driver_mux_selector);
			track_7_3_chanY_n9  <= track_7_3_chanY_n9_driver_mux_fanins(track_7_3_chanY_n9_driver_mux_selector);
			track_7_4_chanX_n0  <= track_7_4_chanX_n0_driver_mux_fanins(track_7_4_chanX_n0_driver_mux_selector);
			track_7_4_chanX_n1  <= track_7_4_chanX_n1_driver_mux_fanins(track_7_4_chanX_n1_driver_mux_selector);
			track_7_4_chanX_n10 <= track_7_4_chanX_n10_driver_mux_fanins(track_7_4_chanX_n10_driver_mux_selector);
			track_7_4_chanX_n11 <= track_7_4_chanX_n11_driver_mux_fanins(track_7_4_chanX_n11_driver_mux_selector);
			track_7_4_chanX_n12 <= track_7_4_chanX_n12_driver_mux_fanins(track_7_4_chanX_n12_driver_mux_selector);
			track_7_4_chanX_n13 <= track_7_4_chanX_n13_driver_mux_fanins(track_7_4_chanX_n13_driver_mux_selector);
			track_7_4_chanX_n14 <= track_7_4_chanX_n14_driver_mux_fanins(track_7_4_chanX_n14_driver_mux_selector);
			track_7_4_chanX_n15 <= track_7_4_chanX_n15_driver_mux_fanins(track_7_4_chanX_n15_driver_mux_selector);
			track_7_4_chanX_n2  <= track_7_4_chanX_n2_driver_mux_fanins(track_7_4_chanX_n2_driver_mux_selector);
			track_7_4_chanX_n3  <= track_7_4_chanX_n3_driver_mux_fanins(track_7_4_chanX_n3_driver_mux_selector);
			track_7_4_chanX_n4  <= track_7_4_chanX_n4_driver_mux_fanins(track_7_4_chanX_n4_driver_mux_selector);
			track_7_4_chanX_n5  <= track_7_4_chanX_n5_driver_mux_fanins(track_7_4_chanX_n5_driver_mux_selector);
			track_7_4_chanX_n6  <= track_7_4_chanX_n6_driver_mux_fanins(track_7_4_chanX_n6_driver_mux_selector);
			track_7_4_chanX_n7  <= track_7_4_chanX_n7_driver_mux_fanins(track_7_4_chanX_n7_driver_mux_selector);
			track_7_4_chanX_n8  <= track_7_4_chanX_n8_driver_mux_fanins(track_7_4_chanX_n8_driver_mux_selector);
			track_7_4_chanX_n9  <= track_7_4_chanX_n9_driver_mux_fanins(track_7_4_chanX_n9_driver_mux_selector);
			track_7_4_chanY_n0  <= track_7_4_chanY_n0_driver_mux_fanins(track_7_4_chanY_n0_driver_mux_selector);
			track_7_4_chanY_n1  <= track_7_4_chanY_n1_driver_mux_fanins(track_7_4_chanY_n1_driver_mux_selector);
			track_7_4_chanY_n10 <= track_7_4_chanY_n10_driver_mux_fanins(track_7_4_chanY_n10_driver_mux_selector);
			track_7_4_chanY_n11 <= track_7_4_chanY_n11_driver_mux_fanins(track_7_4_chanY_n11_driver_mux_selector);
			track_7_4_chanY_n12 <= track_7_4_chanY_n12_driver_mux_fanins(track_7_4_chanY_n12_driver_mux_selector);
			track_7_4_chanY_n13 <= track_7_4_chanY_n13_driver_mux_fanins(track_7_4_chanY_n13_driver_mux_selector);
			track_7_4_chanY_n14 <= track_7_4_chanY_n14_driver_mux_fanins(track_7_4_chanY_n14_driver_mux_selector);
			track_7_4_chanY_n15 <= track_7_4_chanY_n15_driver_mux_fanins(track_7_4_chanY_n15_driver_mux_selector);
			track_7_4_chanY_n2  <= track_7_4_chanY_n2_driver_mux_fanins(track_7_4_chanY_n2_driver_mux_selector);
			track_7_4_chanY_n3  <= track_7_4_chanY_n3_driver_mux_fanins(track_7_4_chanY_n3_driver_mux_selector);
			track_7_4_chanY_n4  <= track_7_4_chanY_n4_driver_mux_fanins(track_7_4_chanY_n4_driver_mux_selector);
			track_7_4_chanY_n5  <= track_7_4_chanY_n5_driver_mux_fanins(track_7_4_chanY_n5_driver_mux_selector);
			track_7_4_chanY_n6  <= track_7_4_chanY_n6_driver_mux_fanins(track_7_4_chanY_n6_driver_mux_selector);
			track_7_4_chanY_n7  <= track_7_4_chanY_n7_driver_mux_fanins(track_7_4_chanY_n7_driver_mux_selector);
			track_7_4_chanY_n8  <= track_7_4_chanY_n8_driver_mux_fanins(track_7_4_chanY_n8_driver_mux_selector);
			track_7_4_chanY_n9  <= track_7_4_chanY_n9_driver_mux_fanins(track_7_4_chanY_n9_driver_mux_selector);
			track_7_5_chanX_n0  <= track_7_5_chanX_n0_driver_mux_fanins(track_7_5_chanX_n0_driver_mux_selector);
			track_7_5_chanX_n1  <= track_7_5_chanX_n1_driver_mux_fanins(track_7_5_chanX_n1_driver_mux_selector);
			track_7_5_chanX_n10 <= track_7_5_chanX_n10_driver_mux_fanins(track_7_5_chanX_n10_driver_mux_selector);
			track_7_5_chanX_n11 <= track_7_5_chanX_n11_driver_mux_fanins(track_7_5_chanX_n11_driver_mux_selector);
			track_7_5_chanX_n12 <= track_7_5_chanX_n12_driver_mux_fanins(track_7_5_chanX_n12_driver_mux_selector);
			track_7_5_chanX_n13 <= track_7_5_chanX_n13_driver_mux_fanins(track_7_5_chanX_n13_driver_mux_selector);
			track_7_5_chanX_n14 <= track_7_5_chanX_n14_driver_mux_fanins(track_7_5_chanX_n14_driver_mux_selector);
			track_7_5_chanX_n15 <= track_7_5_chanX_n15_driver_mux_fanins(track_7_5_chanX_n15_driver_mux_selector);
			track_7_5_chanX_n2  <= track_7_5_chanX_n2_driver_mux_fanins(track_7_5_chanX_n2_driver_mux_selector);
			track_7_5_chanX_n3  <= track_7_5_chanX_n3_driver_mux_fanins(track_7_5_chanX_n3_driver_mux_selector);
			track_7_5_chanX_n4  <= track_7_5_chanX_n4_driver_mux_fanins(track_7_5_chanX_n4_driver_mux_selector);
			track_7_5_chanX_n5  <= track_7_5_chanX_n5_driver_mux_fanins(track_7_5_chanX_n5_driver_mux_selector);
			track_7_5_chanX_n6  <= track_7_5_chanX_n6_driver_mux_fanins(track_7_5_chanX_n6_driver_mux_selector);
			track_7_5_chanX_n7  <= track_7_5_chanX_n7_driver_mux_fanins(track_7_5_chanX_n7_driver_mux_selector);
			track_7_5_chanX_n8  <= track_7_5_chanX_n8_driver_mux_fanins(track_7_5_chanX_n8_driver_mux_selector);
			track_7_5_chanX_n9  <= track_7_5_chanX_n9_driver_mux_fanins(track_7_5_chanX_n9_driver_mux_selector);
			track_7_5_chanY_n0  <= track_7_5_chanY_n0_driver_mux_fanins(track_7_5_chanY_n0_driver_mux_selector);
			track_7_5_chanY_n1  <= track_7_5_chanY_n1_driver_mux_fanins(track_7_5_chanY_n1_driver_mux_selector);
			track_7_5_chanY_n10 <= track_7_5_chanY_n10_driver_mux_fanins(track_7_5_chanY_n10_driver_mux_selector);
			track_7_5_chanY_n11 <= track_7_5_chanY_n11_driver_mux_fanins(track_7_5_chanY_n11_driver_mux_selector);
			track_7_5_chanY_n12 <= track_7_5_chanY_n12_driver_mux_fanins(track_7_5_chanY_n12_driver_mux_selector);
			track_7_5_chanY_n13 <= track_7_5_chanY_n13_driver_mux_fanins(track_7_5_chanY_n13_driver_mux_selector);
			track_7_5_chanY_n14 <= track_7_5_chanY_n14_driver_mux_fanins(track_7_5_chanY_n14_driver_mux_selector);
			track_7_5_chanY_n15 <= track_7_5_chanY_n15_driver_mux_fanins(track_7_5_chanY_n15_driver_mux_selector);
			track_7_5_chanY_n2  <= track_7_5_chanY_n2_driver_mux_fanins(track_7_5_chanY_n2_driver_mux_selector);
			track_7_5_chanY_n3  <= track_7_5_chanY_n3_driver_mux_fanins(track_7_5_chanY_n3_driver_mux_selector);
			track_7_5_chanY_n4  <= track_7_5_chanY_n4_driver_mux_fanins(track_7_5_chanY_n4_driver_mux_selector);
			track_7_5_chanY_n5  <= track_7_5_chanY_n5_driver_mux_fanins(track_7_5_chanY_n5_driver_mux_selector);
			track_7_5_chanY_n6  <= track_7_5_chanY_n6_driver_mux_fanins(track_7_5_chanY_n6_driver_mux_selector);
			track_7_5_chanY_n7  <= track_7_5_chanY_n7_driver_mux_fanins(track_7_5_chanY_n7_driver_mux_selector);
			track_7_5_chanY_n8  <= track_7_5_chanY_n8_driver_mux_fanins(track_7_5_chanY_n8_driver_mux_selector);
			track_7_5_chanY_n9  <= track_7_5_chanY_n9_driver_mux_fanins(track_7_5_chanY_n9_driver_mux_selector);
			track_7_6_chanX_n0  <= track_7_6_chanX_n0_driver_mux_fanins(track_7_6_chanX_n0_driver_mux_selector);
			track_7_6_chanX_n1  <= track_7_6_chanX_n1_driver_mux_fanins(track_7_6_chanX_n1_driver_mux_selector);
			track_7_6_chanX_n10 <= track_7_6_chanX_n10_driver_mux_fanins(track_7_6_chanX_n10_driver_mux_selector);
			track_7_6_chanX_n11 <= track_7_6_chanX_n11_driver_mux_fanins(track_7_6_chanX_n11_driver_mux_selector);
			track_7_6_chanX_n12 <= track_7_6_chanX_n12_driver_mux_fanins(track_7_6_chanX_n12_driver_mux_selector);
			track_7_6_chanX_n13 <= track_7_6_chanX_n13_driver_mux_fanins(track_7_6_chanX_n13_driver_mux_selector);
			track_7_6_chanX_n14 <= track_7_6_chanX_n14_driver_mux_fanins(track_7_6_chanX_n14_driver_mux_selector);
			track_7_6_chanX_n15 <= track_7_6_chanX_n15_driver_mux_fanins(track_7_6_chanX_n15_driver_mux_selector);
			track_7_6_chanX_n2  <= track_7_6_chanX_n2_driver_mux_fanins(track_7_6_chanX_n2_driver_mux_selector);
			track_7_6_chanX_n3  <= track_7_6_chanX_n3_driver_mux_fanins(track_7_6_chanX_n3_driver_mux_selector);
			track_7_6_chanX_n4  <= track_7_6_chanX_n4_driver_mux_fanins(track_7_6_chanX_n4_driver_mux_selector);
			track_7_6_chanX_n5  <= track_7_6_chanX_n5_driver_mux_fanins(track_7_6_chanX_n5_driver_mux_selector);
			track_7_6_chanX_n6  <= track_7_6_chanX_n6_driver_mux_fanins(track_7_6_chanX_n6_driver_mux_selector);
			track_7_6_chanX_n7  <= track_7_6_chanX_n7_driver_mux_fanins(track_7_6_chanX_n7_driver_mux_selector);
			track_7_6_chanX_n8  <= track_7_6_chanX_n8_driver_mux_fanins(track_7_6_chanX_n8_driver_mux_selector);
			track_7_6_chanX_n9  <= track_7_6_chanX_n9_driver_mux_fanins(track_7_6_chanX_n9_driver_mux_selector);
			track_7_6_chanY_n0  <= track_7_6_chanY_n0_driver_mux_fanins(track_7_6_chanY_n0_driver_mux_selector);
			track_7_6_chanY_n1  <= track_7_6_chanY_n1_driver_mux_fanins(track_7_6_chanY_n1_driver_mux_selector);
			track_7_6_chanY_n10 <= track_7_6_chanY_n10_driver_mux_fanins(track_7_6_chanY_n10_driver_mux_selector);
			track_7_6_chanY_n11 <= track_7_6_chanY_n11_driver_mux_fanins(track_7_6_chanY_n11_driver_mux_selector);
			track_7_6_chanY_n12 <= track_7_6_chanY_n12_driver_mux_fanins(track_7_6_chanY_n12_driver_mux_selector);
			track_7_6_chanY_n13 <= track_7_6_chanY_n13_driver_mux_fanins(track_7_6_chanY_n13_driver_mux_selector);
			track_7_6_chanY_n14 <= track_7_6_chanY_n14_driver_mux_fanins(track_7_6_chanY_n14_driver_mux_selector);
			track_7_6_chanY_n15 <= track_7_6_chanY_n15_driver_mux_fanins(track_7_6_chanY_n15_driver_mux_selector);
			track_7_6_chanY_n2  <= track_7_6_chanY_n2_driver_mux_fanins(track_7_6_chanY_n2_driver_mux_selector);
			track_7_6_chanY_n3  <= track_7_6_chanY_n3_driver_mux_fanins(track_7_6_chanY_n3_driver_mux_selector);
			track_7_6_chanY_n4  <= track_7_6_chanY_n4_driver_mux_fanins(track_7_6_chanY_n4_driver_mux_selector);
			track_7_6_chanY_n5  <= track_7_6_chanY_n5_driver_mux_fanins(track_7_6_chanY_n5_driver_mux_selector);
			track_7_6_chanY_n6  <= track_7_6_chanY_n6_driver_mux_fanins(track_7_6_chanY_n6_driver_mux_selector);
			track_7_6_chanY_n7  <= track_7_6_chanY_n7_driver_mux_fanins(track_7_6_chanY_n7_driver_mux_selector);
			track_7_6_chanY_n8  <= track_7_6_chanY_n8_driver_mux_fanins(track_7_6_chanY_n8_driver_mux_selector);
			track_7_6_chanY_n9  <= track_7_6_chanY_n9_driver_mux_fanins(track_7_6_chanY_n9_driver_mux_selector);
			track_8_0_chanX_n0  <= track_8_0_chanX_n0_driver_mux_fanins(track_8_0_chanX_n0_driver_mux_selector);
			track_8_0_chanX_n1  <= track_8_0_chanX_n1_driver_mux_fanins(track_8_0_chanX_n1_driver_mux_selector);
			track_8_0_chanX_n10 <= track_8_0_chanX_n10_driver_mux_fanins(track_8_0_chanX_n10_driver_mux_selector);
			track_8_0_chanX_n11 <= track_8_0_chanX_n11_driver_mux_fanins(track_8_0_chanX_n11_driver_mux_selector);
			track_8_0_chanX_n12 <= track_8_0_chanX_n12_driver_mux_fanins(track_8_0_chanX_n12_driver_mux_selector);
			track_8_0_chanX_n13 <= track_8_0_chanX_n13_driver_mux_fanins(track_8_0_chanX_n13_driver_mux_selector);
			track_8_0_chanX_n14 <= track_8_0_chanX_n14_driver_mux_fanins(track_8_0_chanX_n14_driver_mux_selector);
			track_8_0_chanX_n15 <= track_8_0_chanX_n15_driver_mux_fanins(track_8_0_chanX_n15_driver_mux_selector);
			track_8_0_chanX_n2  <= track_8_0_chanX_n2_driver_mux_fanins(track_8_0_chanX_n2_driver_mux_selector);
			track_8_0_chanX_n3  <= track_8_0_chanX_n3_driver_mux_fanins(track_8_0_chanX_n3_driver_mux_selector);
			track_8_0_chanX_n4  <= track_8_0_chanX_n4_driver_mux_fanins(track_8_0_chanX_n4_driver_mux_selector);
			track_8_0_chanX_n5  <= track_8_0_chanX_n5_driver_mux_fanins(track_8_0_chanX_n5_driver_mux_selector);
			track_8_0_chanX_n6  <= track_8_0_chanX_n6_driver_mux_fanins(track_8_0_chanX_n6_driver_mux_selector);
			track_8_0_chanX_n7  <= track_8_0_chanX_n7_driver_mux_fanins(track_8_0_chanX_n7_driver_mux_selector);
			track_8_0_chanX_n8  <= track_8_0_chanX_n8_driver_mux_fanins(track_8_0_chanX_n8_driver_mux_selector);
			track_8_0_chanX_n9  <= track_8_0_chanX_n9_driver_mux_fanins(track_8_0_chanX_n9_driver_mux_selector);
			track_8_1_chanX_n0  <= track_8_1_chanX_n0_driver_mux_fanins(track_8_1_chanX_n0_driver_mux_selector);
			track_8_1_chanX_n1  <= track_8_1_chanX_n1_driver_mux_fanins(track_8_1_chanX_n1_driver_mux_selector);
			track_8_1_chanX_n10 <= track_8_1_chanX_n10_driver_mux_fanins(track_8_1_chanX_n10_driver_mux_selector);
			track_8_1_chanX_n11 <= track_8_1_chanX_n11_driver_mux_fanins(track_8_1_chanX_n11_driver_mux_selector);
			track_8_1_chanX_n12 <= track_8_1_chanX_n12_driver_mux_fanins(track_8_1_chanX_n12_driver_mux_selector);
			track_8_1_chanX_n13 <= track_8_1_chanX_n13_driver_mux_fanins(track_8_1_chanX_n13_driver_mux_selector);
			track_8_1_chanX_n14 <= track_8_1_chanX_n14_driver_mux_fanins(track_8_1_chanX_n14_driver_mux_selector);
			track_8_1_chanX_n15 <= track_8_1_chanX_n15_driver_mux_fanins(track_8_1_chanX_n15_driver_mux_selector);
			track_8_1_chanX_n2  <= track_8_1_chanX_n2_driver_mux_fanins(track_8_1_chanX_n2_driver_mux_selector);
			track_8_1_chanX_n3  <= track_8_1_chanX_n3_driver_mux_fanins(track_8_1_chanX_n3_driver_mux_selector);
			track_8_1_chanX_n4  <= track_8_1_chanX_n4_driver_mux_fanins(track_8_1_chanX_n4_driver_mux_selector);
			track_8_1_chanX_n5  <= track_8_1_chanX_n5_driver_mux_fanins(track_8_1_chanX_n5_driver_mux_selector);
			track_8_1_chanX_n6  <= track_8_1_chanX_n6_driver_mux_fanins(track_8_1_chanX_n6_driver_mux_selector);
			track_8_1_chanX_n7  <= track_8_1_chanX_n7_driver_mux_fanins(track_8_1_chanX_n7_driver_mux_selector);
			track_8_1_chanX_n8  <= track_8_1_chanX_n8_driver_mux_fanins(track_8_1_chanX_n8_driver_mux_selector);
			track_8_1_chanX_n9  <= track_8_1_chanX_n9_driver_mux_fanins(track_8_1_chanX_n9_driver_mux_selector);
			track_8_1_chanY_n0  <= track_8_1_chanY_n0_driver_mux_fanins(track_8_1_chanY_n0_driver_mux_selector);
			track_8_1_chanY_n1  <= track_8_1_chanY_n1_driver_mux_fanins(track_8_1_chanY_n1_driver_mux_selector);
			track_8_1_chanY_n10 <= track_8_1_chanY_n10_driver_mux_fanins(track_8_1_chanY_n10_driver_mux_selector);
			track_8_1_chanY_n11 <= track_8_1_chanY_n11_driver_mux_fanins(track_8_1_chanY_n11_driver_mux_selector);
			track_8_1_chanY_n12 <= track_8_1_chanY_n12_driver_mux_fanins(track_8_1_chanY_n12_driver_mux_selector);
			track_8_1_chanY_n13 <= track_8_1_chanY_n13_driver_mux_fanins(track_8_1_chanY_n13_driver_mux_selector);
			track_8_1_chanY_n14 <= track_8_1_chanY_n14_driver_mux_fanins(track_8_1_chanY_n14_driver_mux_selector);
			track_8_1_chanY_n15 <= track_8_1_chanY_n15_driver_mux_fanins(track_8_1_chanY_n15_driver_mux_selector);
			track_8_1_chanY_n2  <= track_8_1_chanY_n2_driver_mux_fanins(track_8_1_chanY_n2_driver_mux_selector);
			track_8_1_chanY_n3  <= track_8_1_chanY_n3_driver_mux_fanins(track_8_1_chanY_n3_driver_mux_selector);
			track_8_1_chanY_n4  <= track_8_1_chanY_n4_driver_mux_fanins(track_8_1_chanY_n4_driver_mux_selector);
			track_8_1_chanY_n5  <= track_8_1_chanY_n5_driver_mux_fanins(track_8_1_chanY_n5_driver_mux_selector);
			track_8_1_chanY_n6  <= track_8_1_chanY_n6_driver_mux_fanins(track_8_1_chanY_n6_driver_mux_selector);
			track_8_1_chanY_n7  <= track_8_1_chanY_n7_driver_mux_fanins(track_8_1_chanY_n7_driver_mux_selector);
			track_8_1_chanY_n8  <= track_8_1_chanY_n8_driver_mux_fanins(track_8_1_chanY_n8_driver_mux_selector);
			track_8_1_chanY_n9  <= track_8_1_chanY_n9_driver_mux_fanins(track_8_1_chanY_n9_driver_mux_selector);
			track_8_2_chanX_n0  <= track_8_2_chanX_n0_driver_mux_fanins(track_8_2_chanX_n0_driver_mux_selector);
			track_8_2_chanX_n1  <= track_8_2_chanX_n1_driver_mux_fanins(track_8_2_chanX_n1_driver_mux_selector);
			track_8_2_chanX_n10 <= track_8_2_chanX_n10_driver_mux_fanins(track_8_2_chanX_n10_driver_mux_selector);
			track_8_2_chanX_n11 <= track_8_2_chanX_n11_driver_mux_fanins(track_8_2_chanX_n11_driver_mux_selector);
			track_8_2_chanX_n12 <= track_8_2_chanX_n12_driver_mux_fanins(track_8_2_chanX_n12_driver_mux_selector);
			track_8_2_chanX_n13 <= track_8_2_chanX_n13_driver_mux_fanins(track_8_2_chanX_n13_driver_mux_selector);
			track_8_2_chanX_n14 <= track_8_2_chanX_n14_driver_mux_fanins(track_8_2_chanX_n14_driver_mux_selector);
			track_8_2_chanX_n15 <= track_8_2_chanX_n15_driver_mux_fanins(track_8_2_chanX_n15_driver_mux_selector);
			track_8_2_chanX_n2  <= track_8_2_chanX_n2_driver_mux_fanins(track_8_2_chanX_n2_driver_mux_selector);
			track_8_2_chanX_n3  <= track_8_2_chanX_n3_driver_mux_fanins(track_8_2_chanX_n3_driver_mux_selector);
			track_8_2_chanX_n4  <= track_8_2_chanX_n4_driver_mux_fanins(track_8_2_chanX_n4_driver_mux_selector);
			track_8_2_chanX_n5  <= track_8_2_chanX_n5_driver_mux_fanins(track_8_2_chanX_n5_driver_mux_selector);
			track_8_2_chanX_n6  <= track_8_2_chanX_n6_driver_mux_fanins(track_8_2_chanX_n6_driver_mux_selector);
			track_8_2_chanX_n7  <= track_8_2_chanX_n7_driver_mux_fanins(track_8_2_chanX_n7_driver_mux_selector);
			track_8_2_chanX_n8  <= track_8_2_chanX_n8_driver_mux_fanins(track_8_2_chanX_n8_driver_mux_selector);
			track_8_2_chanX_n9  <= track_8_2_chanX_n9_driver_mux_fanins(track_8_2_chanX_n9_driver_mux_selector);
			track_8_2_chanY_n0  <= track_8_2_chanY_n0_driver_mux_fanins(track_8_2_chanY_n0_driver_mux_selector);
			track_8_2_chanY_n1  <= track_8_2_chanY_n1_driver_mux_fanins(track_8_2_chanY_n1_driver_mux_selector);
			track_8_2_chanY_n10 <= track_8_2_chanY_n10_driver_mux_fanins(track_8_2_chanY_n10_driver_mux_selector);
			track_8_2_chanY_n11 <= track_8_2_chanY_n11_driver_mux_fanins(track_8_2_chanY_n11_driver_mux_selector);
			track_8_2_chanY_n12 <= track_8_2_chanY_n12_driver_mux_fanins(track_8_2_chanY_n12_driver_mux_selector);
			track_8_2_chanY_n13 <= track_8_2_chanY_n13_driver_mux_fanins(track_8_2_chanY_n13_driver_mux_selector);
			track_8_2_chanY_n14 <= track_8_2_chanY_n14_driver_mux_fanins(track_8_2_chanY_n14_driver_mux_selector);
			track_8_2_chanY_n15 <= track_8_2_chanY_n15_driver_mux_fanins(track_8_2_chanY_n15_driver_mux_selector);
			track_8_2_chanY_n2  <= track_8_2_chanY_n2_driver_mux_fanins(track_8_2_chanY_n2_driver_mux_selector);
			track_8_2_chanY_n3  <= track_8_2_chanY_n3_driver_mux_fanins(track_8_2_chanY_n3_driver_mux_selector);
			track_8_2_chanY_n4  <= track_8_2_chanY_n4_driver_mux_fanins(track_8_2_chanY_n4_driver_mux_selector);
			track_8_2_chanY_n5  <= track_8_2_chanY_n5_driver_mux_fanins(track_8_2_chanY_n5_driver_mux_selector);
			track_8_2_chanY_n6  <= track_8_2_chanY_n6_driver_mux_fanins(track_8_2_chanY_n6_driver_mux_selector);
			track_8_2_chanY_n7  <= track_8_2_chanY_n7_driver_mux_fanins(track_8_2_chanY_n7_driver_mux_selector);
			track_8_2_chanY_n8  <= track_8_2_chanY_n8_driver_mux_fanins(track_8_2_chanY_n8_driver_mux_selector);
			track_8_2_chanY_n9  <= track_8_2_chanY_n9_driver_mux_fanins(track_8_2_chanY_n9_driver_mux_selector);
			track_8_3_chanX_n0  <= track_8_3_chanX_n0_driver_mux_fanins(track_8_3_chanX_n0_driver_mux_selector);
			track_8_3_chanX_n1  <= track_8_3_chanX_n1_driver_mux_fanins(track_8_3_chanX_n1_driver_mux_selector);
			track_8_3_chanX_n10 <= track_8_3_chanX_n10_driver_mux_fanins(track_8_3_chanX_n10_driver_mux_selector);
			track_8_3_chanX_n11 <= track_8_3_chanX_n11_driver_mux_fanins(track_8_3_chanX_n11_driver_mux_selector);
			track_8_3_chanX_n12 <= track_8_3_chanX_n12_driver_mux_fanins(track_8_3_chanX_n12_driver_mux_selector);
			track_8_3_chanX_n13 <= track_8_3_chanX_n13_driver_mux_fanins(track_8_3_chanX_n13_driver_mux_selector);
			track_8_3_chanX_n14 <= track_8_3_chanX_n14_driver_mux_fanins(track_8_3_chanX_n14_driver_mux_selector);
			track_8_3_chanX_n15 <= track_8_3_chanX_n15_driver_mux_fanins(track_8_3_chanX_n15_driver_mux_selector);
			track_8_3_chanX_n2  <= track_8_3_chanX_n2_driver_mux_fanins(track_8_3_chanX_n2_driver_mux_selector);
			track_8_3_chanX_n3  <= track_8_3_chanX_n3_driver_mux_fanins(track_8_3_chanX_n3_driver_mux_selector);
			track_8_3_chanX_n4  <= track_8_3_chanX_n4_driver_mux_fanins(track_8_3_chanX_n4_driver_mux_selector);
			track_8_3_chanX_n5  <= track_8_3_chanX_n5_driver_mux_fanins(track_8_3_chanX_n5_driver_mux_selector);
			track_8_3_chanX_n6  <= track_8_3_chanX_n6_driver_mux_fanins(track_8_3_chanX_n6_driver_mux_selector);
			track_8_3_chanX_n7  <= track_8_3_chanX_n7_driver_mux_fanins(track_8_3_chanX_n7_driver_mux_selector);
			track_8_3_chanX_n8  <= track_8_3_chanX_n8_driver_mux_fanins(track_8_3_chanX_n8_driver_mux_selector);
			track_8_3_chanX_n9  <= track_8_3_chanX_n9_driver_mux_fanins(track_8_3_chanX_n9_driver_mux_selector);
			track_8_3_chanY_n0  <= track_8_3_chanY_n0_driver_mux_fanins(track_8_3_chanY_n0_driver_mux_selector);
			track_8_3_chanY_n1  <= track_8_3_chanY_n1_driver_mux_fanins(track_8_3_chanY_n1_driver_mux_selector);
			track_8_3_chanY_n10 <= track_8_3_chanY_n10_driver_mux_fanins(track_8_3_chanY_n10_driver_mux_selector);
			track_8_3_chanY_n11 <= track_8_3_chanY_n11_driver_mux_fanins(track_8_3_chanY_n11_driver_mux_selector);
			track_8_3_chanY_n12 <= track_8_3_chanY_n12_driver_mux_fanins(track_8_3_chanY_n12_driver_mux_selector);
			track_8_3_chanY_n13 <= track_8_3_chanY_n13_driver_mux_fanins(track_8_3_chanY_n13_driver_mux_selector);
			track_8_3_chanY_n14 <= track_8_3_chanY_n14_driver_mux_fanins(track_8_3_chanY_n14_driver_mux_selector);
			track_8_3_chanY_n15 <= track_8_3_chanY_n15_driver_mux_fanins(track_8_3_chanY_n15_driver_mux_selector);
			track_8_3_chanY_n2  <= track_8_3_chanY_n2_driver_mux_fanins(track_8_3_chanY_n2_driver_mux_selector);
			track_8_3_chanY_n3  <= track_8_3_chanY_n3_driver_mux_fanins(track_8_3_chanY_n3_driver_mux_selector);
			track_8_3_chanY_n4  <= track_8_3_chanY_n4_driver_mux_fanins(track_8_3_chanY_n4_driver_mux_selector);
			track_8_3_chanY_n5  <= track_8_3_chanY_n5_driver_mux_fanins(track_8_3_chanY_n5_driver_mux_selector);
			track_8_3_chanY_n6  <= track_8_3_chanY_n6_driver_mux_fanins(track_8_3_chanY_n6_driver_mux_selector);
			track_8_3_chanY_n7  <= track_8_3_chanY_n7_driver_mux_fanins(track_8_3_chanY_n7_driver_mux_selector);
			track_8_3_chanY_n8  <= track_8_3_chanY_n8_driver_mux_fanins(track_8_3_chanY_n8_driver_mux_selector);
			track_8_3_chanY_n9  <= track_8_3_chanY_n9_driver_mux_fanins(track_8_3_chanY_n9_driver_mux_selector);
			track_8_4_chanX_n0  <= track_8_4_chanX_n0_driver_mux_fanins(track_8_4_chanX_n0_driver_mux_selector);
			track_8_4_chanX_n1  <= track_8_4_chanX_n1_driver_mux_fanins(track_8_4_chanX_n1_driver_mux_selector);
			track_8_4_chanX_n10 <= track_8_4_chanX_n10_driver_mux_fanins(track_8_4_chanX_n10_driver_mux_selector);
			track_8_4_chanX_n11 <= track_8_4_chanX_n11_driver_mux_fanins(track_8_4_chanX_n11_driver_mux_selector);
			track_8_4_chanX_n12 <= track_8_4_chanX_n12_driver_mux_fanins(track_8_4_chanX_n12_driver_mux_selector);
			track_8_4_chanX_n13 <= track_8_4_chanX_n13_driver_mux_fanins(track_8_4_chanX_n13_driver_mux_selector);
			track_8_4_chanX_n14 <= track_8_4_chanX_n14_driver_mux_fanins(track_8_4_chanX_n14_driver_mux_selector);
			track_8_4_chanX_n15 <= track_8_4_chanX_n15_driver_mux_fanins(track_8_4_chanX_n15_driver_mux_selector);
			track_8_4_chanX_n2  <= track_8_4_chanX_n2_driver_mux_fanins(track_8_4_chanX_n2_driver_mux_selector);
			track_8_4_chanX_n3  <= track_8_4_chanX_n3_driver_mux_fanins(track_8_4_chanX_n3_driver_mux_selector);
			track_8_4_chanX_n4  <= track_8_4_chanX_n4_driver_mux_fanins(track_8_4_chanX_n4_driver_mux_selector);
			track_8_4_chanX_n5  <= track_8_4_chanX_n5_driver_mux_fanins(track_8_4_chanX_n5_driver_mux_selector);
			track_8_4_chanX_n6  <= track_8_4_chanX_n6_driver_mux_fanins(track_8_4_chanX_n6_driver_mux_selector);
			track_8_4_chanX_n7  <= track_8_4_chanX_n7_driver_mux_fanins(track_8_4_chanX_n7_driver_mux_selector);
			track_8_4_chanX_n8  <= track_8_4_chanX_n8_driver_mux_fanins(track_8_4_chanX_n8_driver_mux_selector);
			track_8_4_chanX_n9  <= track_8_4_chanX_n9_driver_mux_fanins(track_8_4_chanX_n9_driver_mux_selector);
			track_8_4_chanY_n0  <= track_8_4_chanY_n0_driver_mux_fanins(track_8_4_chanY_n0_driver_mux_selector);
			track_8_4_chanY_n1  <= track_8_4_chanY_n1_driver_mux_fanins(track_8_4_chanY_n1_driver_mux_selector);
			track_8_4_chanY_n10 <= track_8_4_chanY_n10_driver_mux_fanins(track_8_4_chanY_n10_driver_mux_selector);
			track_8_4_chanY_n11 <= track_8_4_chanY_n11_driver_mux_fanins(track_8_4_chanY_n11_driver_mux_selector);
			track_8_4_chanY_n12 <= track_8_4_chanY_n12_driver_mux_fanins(track_8_4_chanY_n12_driver_mux_selector);
			track_8_4_chanY_n13 <= track_8_4_chanY_n13_driver_mux_fanins(track_8_4_chanY_n13_driver_mux_selector);
			track_8_4_chanY_n14 <= track_8_4_chanY_n14_driver_mux_fanins(track_8_4_chanY_n14_driver_mux_selector);
			track_8_4_chanY_n15 <= track_8_4_chanY_n15_driver_mux_fanins(track_8_4_chanY_n15_driver_mux_selector);
			track_8_4_chanY_n2  <= track_8_4_chanY_n2_driver_mux_fanins(track_8_4_chanY_n2_driver_mux_selector);
			track_8_4_chanY_n3  <= track_8_4_chanY_n3_driver_mux_fanins(track_8_4_chanY_n3_driver_mux_selector);
			track_8_4_chanY_n4  <= track_8_4_chanY_n4_driver_mux_fanins(track_8_4_chanY_n4_driver_mux_selector);
			track_8_4_chanY_n5  <= track_8_4_chanY_n5_driver_mux_fanins(track_8_4_chanY_n5_driver_mux_selector);
			track_8_4_chanY_n6  <= track_8_4_chanY_n6_driver_mux_fanins(track_8_4_chanY_n6_driver_mux_selector);
			track_8_4_chanY_n7  <= track_8_4_chanY_n7_driver_mux_fanins(track_8_4_chanY_n7_driver_mux_selector);
			track_8_4_chanY_n8  <= track_8_4_chanY_n8_driver_mux_fanins(track_8_4_chanY_n8_driver_mux_selector);
			track_8_4_chanY_n9  <= track_8_4_chanY_n9_driver_mux_fanins(track_8_4_chanY_n9_driver_mux_selector);
			track_8_5_chanX_n0  <= track_8_5_chanX_n0_driver_mux_fanins(track_8_5_chanX_n0_driver_mux_selector);
			track_8_5_chanX_n1  <= track_8_5_chanX_n1_driver_mux_fanins(track_8_5_chanX_n1_driver_mux_selector);
			track_8_5_chanX_n10 <= track_8_5_chanX_n10_driver_mux_fanins(track_8_5_chanX_n10_driver_mux_selector);
			track_8_5_chanX_n11 <= track_8_5_chanX_n11_driver_mux_fanins(track_8_5_chanX_n11_driver_mux_selector);
			track_8_5_chanX_n12 <= track_8_5_chanX_n12_driver_mux_fanins(track_8_5_chanX_n12_driver_mux_selector);
			track_8_5_chanX_n13 <= track_8_5_chanX_n13_driver_mux_fanins(track_8_5_chanX_n13_driver_mux_selector);
			track_8_5_chanX_n14 <= track_8_5_chanX_n14_driver_mux_fanins(track_8_5_chanX_n14_driver_mux_selector);
			track_8_5_chanX_n15 <= track_8_5_chanX_n15_driver_mux_fanins(track_8_5_chanX_n15_driver_mux_selector);
			track_8_5_chanX_n2  <= track_8_5_chanX_n2_driver_mux_fanins(track_8_5_chanX_n2_driver_mux_selector);
			track_8_5_chanX_n3  <= track_8_5_chanX_n3_driver_mux_fanins(track_8_5_chanX_n3_driver_mux_selector);
			track_8_5_chanX_n4  <= track_8_5_chanX_n4_driver_mux_fanins(track_8_5_chanX_n4_driver_mux_selector);
			track_8_5_chanX_n5  <= track_8_5_chanX_n5_driver_mux_fanins(track_8_5_chanX_n5_driver_mux_selector);
			track_8_5_chanX_n6  <= track_8_5_chanX_n6_driver_mux_fanins(track_8_5_chanX_n6_driver_mux_selector);
			track_8_5_chanX_n7  <= track_8_5_chanX_n7_driver_mux_fanins(track_8_5_chanX_n7_driver_mux_selector);
			track_8_5_chanX_n8  <= track_8_5_chanX_n8_driver_mux_fanins(track_8_5_chanX_n8_driver_mux_selector);
			track_8_5_chanX_n9  <= track_8_5_chanX_n9_driver_mux_fanins(track_8_5_chanX_n9_driver_mux_selector);
			track_8_5_chanY_n0  <= track_8_5_chanY_n0_driver_mux_fanins(track_8_5_chanY_n0_driver_mux_selector);
			track_8_5_chanY_n1  <= track_8_5_chanY_n1_driver_mux_fanins(track_8_5_chanY_n1_driver_mux_selector);
			track_8_5_chanY_n10 <= track_8_5_chanY_n10_driver_mux_fanins(track_8_5_chanY_n10_driver_mux_selector);
			track_8_5_chanY_n11 <= track_8_5_chanY_n11_driver_mux_fanins(track_8_5_chanY_n11_driver_mux_selector);
			track_8_5_chanY_n12 <= track_8_5_chanY_n12_driver_mux_fanins(track_8_5_chanY_n12_driver_mux_selector);
			track_8_5_chanY_n13 <= track_8_5_chanY_n13_driver_mux_fanins(track_8_5_chanY_n13_driver_mux_selector);
			track_8_5_chanY_n14 <= track_8_5_chanY_n14_driver_mux_fanins(track_8_5_chanY_n14_driver_mux_selector);
			track_8_5_chanY_n15 <= track_8_5_chanY_n15_driver_mux_fanins(track_8_5_chanY_n15_driver_mux_selector);
			track_8_5_chanY_n2  <= track_8_5_chanY_n2_driver_mux_fanins(track_8_5_chanY_n2_driver_mux_selector);
			track_8_5_chanY_n3  <= track_8_5_chanY_n3_driver_mux_fanins(track_8_5_chanY_n3_driver_mux_selector);
			track_8_5_chanY_n4  <= track_8_5_chanY_n4_driver_mux_fanins(track_8_5_chanY_n4_driver_mux_selector);
			track_8_5_chanY_n5  <= track_8_5_chanY_n5_driver_mux_fanins(track_8_5_chanY_n5_driver_mux_selector);
			track_8_5_chanY_n6  <= track_8_5_chanY_n6_driver_mux_fanins(track_8_5_chanY_n6_driver_mux_selector);
			track_8_5_chanY_n7  <= track_8_5_chanY_n7_driver_mux_fanins(track_8_5_chanY_n7_driver_mux_selector);
			track_8_5_chanY_n8  <= track_8_5_chanY_n8_driver_mux_fanins(track_8_5_chanY_n8_driver_mux_selector);
			track_8_5_chanY_n9  <= track_8_5_chanY_n9_driver_mux_fanins(track_8_5_chanY_n9_driver_mux_selector);
			track_8_6_chanX_n0  <= track_8_6_chanX_n0_driver_mux_fanins(track_8_6_chanX_n0_driver_mux_selector);
			track_8_6_chanX_n1  <= track_8_6_chanX_n1_driver_mux_fanins(track_8_6_chanX_n1_driver_mux_selector);
			track_8_6_chanX_n10 <= track_8_6_chanX_n10_driver_mux_fanins(track_8_6_chanX_n10_driver_mux_selector);
			track_8_6_chanX_n11 <= track_8_6_chanX_n11_driver_mux_fanins(track_8_6_chanX_n11_driver_mux_selector);
			track_8_6_chanX_n12 <= track_8_6_chanX_n12_driver_mux_fanins(track_8_6_chanX_n12_driver_mux_selector);
			track_8_6_chanX_n13 <= track_8_6_chanX_n13_driver_mux_fanins(track_8_6_chanX_n13_driver_mux_selector);
			track_8_6_chanX_n14 <= track_8_6_chanX_n14_driver_mux_fanins(track_8_6_chanX_n14_driver_mux_selector);
			track_8_6_chanX_n15 <= track_8_6_chanX_n15_driver_mux_fanins(track_8_6_chanX_n15_driver_mux_selector);
			track_8_6_chanX_n2  <= track_8_6_chanX_n2_driver_mux_fanins(track_8_6_chanX_n2_driver_mux_selector);
			track_8_6_chanX_n3  <= track_8_6_chanX_n3_driver_mux_fanins(track_8_6_chanX_n3_driver_mux_selector);
			track_8_6_chanX_n4  <= track_8_6_chanX_n4_driver_mux_fanins(track_8_6_chanX_n4_driver_mux_selector);
			track_8_6_chanX_n5  <= track_8_6_chanX_n5_driver_mux_fanins(track_8_6_chanX_n5_driver_mux_selector);
			track_8_6_chanX_n6  <= track_8_6_chanX_n6_driver_mux_fanins(track_8_6_chanX_n6_driver_mux_selector);
			track_8_6_chanX_n7  <= track_8_6_chanX_n7_driver_mux_fanins(track_8_6_chanX_n7_driver_mux_selector);
			track_8_6_chanX_n8  <= track_8_6_chanX_n8_driver_mux_fanins(track_8_6_chanX_n8_driver_mux_selector);
			track_8_6_chanX_n9  <= track_8_6_chanX_n9_driver_mux_fanins(track_8_6_chanX_n9_driver_mux_selector);
			track_8_6_chanY_n0  <= track_8_6_chanY_n0_driver_mux_fanins(track_8_6_chanY_n0_driver_mux_selector);
			track_8_6_chanY_n1  <= track_8_6_chanY_n1_driver_mux_fanins(track_8_6_chanY_n1_driver_mux_selector);
			track_8_6_chanY_n10 <= track_8_6_chanY_n10_driver_mux_fanins(track_8_6_chanY_n10_driver_mux_selector);
			track_8_6_chanY_n11 <= track_8_6_chanY_n11_driver_mux_fanins(track_8_6_chanY_n11_driver_mux_selector);
			track_8_6_chanY_n12 <= track_8_6_chanY_n12_driver_mux_fanins(track_8_6_chanY_n12_driver_mux_selector);
			track_8_6_chanY_n13 <= track_8_6_chanY_n13_driver_mux_fanins(track_8_6_chanY_n13_driver_mux_selector);
			track_8_6_chanY_n14 <= track_8_6_chanY_n14_driver_mux_fanins(track_8_6_chanY_n14_driver_mux_selector);
			track_8_6_chanY_n15 <= track_8_6_chanY_n15_driver_mux_fanins(track_8_6_chanY_n15_driver_mux_selector);
			track_8_6_chanY_n2  <= track_8_6_chanY_n2_driver_mux_fanins(track_8_6_chanY_n2_driver_mux_selector);
			track_8_6_chanY_n3  <= track_8_6_chanY_n3_driver_mux_fanins(track_8_6_chanY_n3_driver_mux_selector);
			track_8_6_chanY_n4  <= track_8_6_chanY_n4_driver_mux_fanins(track_8_6_chanY_n4_driver_mux_selector);
			track_8_6_chanY_n5  <= track_8_6_chanY_n5_driver_mux_fanins(track_8_6_chanY_n5_driver_mux_selector);
			track_8_6_chanY_n6  <= track_8_6_chanY_n6_driver_mux_fanins(track_8_6_chanY_n6_driver_mux_selector);
			track_8_6_chanY_n7  <= track_8_6_chanY_n7_driver_mux_fanins(track_8_6_chanY_n7_driver_mux_selector);
			track_8_6_chanY_n8  <= track_8_6_chanY_n8_driver_mux_fanins(track_8_6_chanY_n8_driver_mux_selector);
			track_8_6_chanY_n9  <= track_8_6_chanY_n9_driver_mux_fanins(track_8_6_chanY_n9_driver_mux_selector);
		end if;
	end process;

	-- vFPGA output pads --
	outputs(55) <= IO_0_1_IN_pin_0;
	outputs(54) <= IO_0_1_IN_pin_1;
	outputs(53) <= IO_0_2_IN_pin_0;
	outputs(52) <= IO_0_2_IN_pin_1;
	outputs(51) <= IO_0_3_IN_pin_0;
	outputs(50) <= IO_0_3_IN_pin_1;
	outputs(49) <= IO_0_4_IN_pin_0;
	outputs(48) <= IO_0_4_IN_pin_1;
	outputs(47) <= IO_0_5_IN_pin_0;
	outputs(46) <= IO_0_5_IN_pin_1;
	outputs(45) <= IO_0_6_IN_pin_0;
	outputs(44) <= IO_0_6_IN_pin_1;
	outputs(43) <= IO_1_7_IN_pin_0;
	outputs(42) <= IO_1_7_IN_pin_1;
	outputs(41) <= IO_2_7_IN_pin_0;
	outputs(40) <= IO_2_7_IN_pin_1;
	outputs(39) <= IO_3_7_IN_pin_0;
	outputs(38) <= IO_3_7_IN_pin_1;
	outputs(37) <= IO_4_7_IN_pin_0;
	outputs(36) <= IO_4_7_IN_pin_1;
	outputs(35) <= IO_5_7_IN_pin_0;
	outputs(34) <= IO_5_7_IN_pin_1;
	outputs(33) <= IO_6_7_IN_pin_0;
	outputs(32) <= IO_6_7_IN_pin_1;
	outputs(31) <= IO_7_7_IN_pin_0;
	outputs(30) <= IO_7_7_IN_pin_1;
	outputs(29) <= IO_8_7_IN_pin_0;
	outputs(28) <= IO_8_7_IN_pin_1;
	outputs(27) <= IO_9_6_IN_pin_1;
	outputs(26) <= IO_9_6_IN_pin_0;
	outputs(25) <= IO_9_5_IN_pin_1;
	outputs(24) <= IO_9_5_IN_pin_0;
	outputs(23) <= IO_9_4_IN_pin_1;
	outputs(22) <= IO_9_4_IN_pin_0;
	outputs(21) <= IO_9_3_IN_pin_1;
	outputs(20) <= IO_9_3_IN_pin_0;
	outputs(19) <= IO_9_2_IN_pin_1;
	outputs(18) <= IO_9_2_IN_pin_0;
	outputs(17) <= IO_9_1_IN_pin_1;
	outputs(16) <= IO_9_1_IN_pin_0;
	outputs(15) <= IO_8_0_IN_pin_1;
	outputs(14) <= IO_8_0_IN_pin_0;
	outputs(13) <= IO_7_0_IN_pin_1;
	outputs(12) <= IO_7_0_IN_pin_0;
	outputs(11) <= IO_6_0_IN_pin_1;
	outputs(10) <= IO_6_0_IN_pin_0;
	outputs( 9) <= IO_5_0_IN_pin_1;
	outputs( 8) <= IO_5_0_IN_pin_0;
	outputs( 7) <= IO_4_0_IN_pin_1;
	outputs( 6) <= IO_4_0_IN_pin_0;
	outputs( 5) <= IO_3_0_IN_pin_1;
	outputs( 4) <= IO_3_0_IN_pin_0;
	outputs( 3) <= IO_2_0_IN_pin_1;
	outputs( 2) <= IO_2_0_IN_pin_0;
	outputs( 1) <= IO_1_0_IN_pin_1;
	outputs( 0) <= IO_1_0_IN_pin_0;

	-- vFPGA input pads --
	IO_0_1_OUT_pin_0 <= inputs(55);
	IO_0_1_OUT_pin_1 <= inputs(54);
	IO_0_2_OUT_pin_0 <= inputs(53);
	IO_0_2_OUT_pin_1 <= inputs(52);
	IO_0_3_OUT_pin_0 <= inputs(51);
	IO_0_3_OUT_pin_1 <= inputs(50);
	IO_0_4_OUT_pin_0 <= inputs(49);
	IO_0_4_OUT_pin_1 <= inputs(48);
	IO_0_5_OUT_pin_0 <= inputs(47);
	IO_0_5_OUT_pin_1 <= inputs(46);
	IO_0_6_OUT_pin_0 <= inputs(45);
	IO_0_6_OUT_pin_1 <= inputs(44);
	IO_1_7_OUT_pin_0 <= inputs(43);
	IO_1_7_OUT_pin_1 <= inputs(42);
	IO_2_7_OUT_pin_0 <= inputs(41);
	IO_2_7_OUT_pin_1 <= inputs(40);
	IO_3_7_OUT_pin_0 <= inputs(39);
	IO_3_7_OUT_pin_1 <= inputs(38);
	IO_4_7_OUT_pin_0 <= inputs(37);
	IO_4_7_OUT_pin_1 <= inputs(36);
	IO_5_7_OUT_pin_0 <= inputs(35);
	IO_5_7_OUT_pin_1 <= inputs(34);
	IO_6_7_OUT_pin_0 <= inputs(33);
	IO_6_7_OUT_pin_1 <= inputs(32);
	IO_7_7_OUT_pin_0 <= inputs(31);
	IO_7_7_OUT_pin_1 <= inputs(30);
	IO_8_7_OUT_pin_0 <= inputs(29);
	IO_8_7_OUT_pin_1 <= inputs(28);
	IO_9_6_OUT_pin_1 <= inputs(27);
	IO_9_6_OUT_pin_0 <= inputs(26);
	IO_9_5_OUT_pin_1 <= inputs(25);
	IO_9_5_OUT_pin_0 <= inputs(24);
	IO_9_4_OUT_pin_1 <= inputs(23);
	IO_9_4_OUT_pin_0 <= inputs(22);
	IO_9_3_OUT_pin_1 <= inputs(21);
	IO_9_3_OUT_pin_0 <= inputs(20);
	IO_9_2_OUT_pin_1 <= inputs(19);
	IO_9_2_OUT_pin_0 <= inputs(18);
	IO_9_1_OUT_pin_1 <= inputs(17);
	IO_9_1_OUT_pin_0 <= inputs(16);
	IO_8_0_OUT_pin_1 <= inputs(15);
	IO_8_0_OUT_pin_0 <= inputs(14);
	IO_7_0_OUT_pin_1 <= inputs(13);
	IO_7_0_OUT_pin_0 <= inputs(12);
	IO_6_0_OUT_pin_1 <= inputs(11);
	IO_6_0_OUT_pin_0 <= inputs(10);
	IO_5_0_OUT_pin_1 <= inputs( 9);
	IO_5_0_OUT_pin_0 <= inputs( 8);
	IO_4_0_OUT_pin_1 <= inputs( 7);
	IO_4_0_OUT_pin_0 <= inputs( 6);
	IO_3_0_OUT_pin_1 <= inputs( 5);
	IO_3_0_OUT_pin_0 <= inputs( 4);
	IO_2_0_OUT_pin_1 <= inputs( 3);
	IO_2_0_OUT_pin_0 <= inputs( 2);
	IO_1_0_OUT_pin_1 <= inputs( 1);
	IO_1_0_OUT_pin_0 <= inputs( 0);

	-- CLB inputs --
	CLB_1_1_inputs <= CLB_1_1_IN_pin_9 & CLB_1_1_IN_pin_8 & CLB_1_1_IN_pin_7 & CLB_1_1_IN_pin_6 & CLB_1_1_IN_pin_5 & CLB_1_1_IN_pin_4 & CLB_1_1_IN_pin_3 & CLB_1_1_IN_pin_2 & CLB_1_1_IN_pin_1 & CLB_1_1_IN_pin_0;
	CLB_1_2_inputs <= CLB_1_2_IN_pin_9 & CLB_1_2_IN_pin_8 & CLB_1_2_IN_pin_7 & CLB_1_2_IN_pin_6 & CLB_1_2_IN_pin_5 & CLB_1_2_IN_pin_4 & CLB_1_2_IN_pin_3 & CLB_1_2_IN_pin_2 & CLB_1_2_IN_pin_1 & CLB_1_2_IN_pin_0;
	CLB_1_3_inputs <= CLB_1_3_IN_pin_9 & CLB_1_3_IN_pin_8 & CLB_1_3_IN_pin_7 & CLB_1_3_IN_pin_6 & CLB_1_3_IN_pin_5 & CLB_1_3_IN_pin_4 & CLB_1_3_IN_pin_3 & CLB_1_3_IN_pin_2 & CLB_1_3_IN_pin_1 & CLB_1_3_IN_pin_0;
	CLB_1_4_inputs <= CLB_1_4_IN_pin_9 & CLB_1_4_IN_pin_8 & CLB_1_4_IN_pin_7 & CLB_1_4_IN_pin_6 & CLB_1_4_IN_pin_5 & CLB_1_4_IN_pin_4 & CLB_1_4_IN_pin_3 & CLB_1_4_IN_pin_2 & CLB_1_4_IN_pin_1 & CLB_1_4_IN_pin_0;
	CLB_1_5_inputs <= CLB_1_5_IN_pin_9 & CLB_1_5_IN_pin_8 & CLB_1_5_IN_pin_7 & CLB_1_5_IN_pin_6 & CLB_1_5_IN_pin_5 & CLB_1_5_IN_pin_4 & CLB_1_5_IN_pin_3 & CLB_1_5_IN_pin_2 & CLB_1_5_IN_pin_1 & CLB_1_5_IN_pin_0;
	CLB_1_6_inputs <= CLB_1_6_IN_pin_9 & CLB_1_6_IN_pin_8 & CLB_1_6_IN_pin_7 & CLB_1_6_IN_pin_6 & CLB_1_6_IN_pin_5 & CLB_1_6_IN_pin_4 & CLB_1_6_IN_pin_3 & CLB_1_6_IN_pin_2 & CLB_1_6_IN_pin_1 & CLB_1_6_IN_pin_0;
	CLB_2_1_inputs <= CLB_2_1_IN_pin_9 & CLB_2_1_IN_pin_8 & CLB_2_1_IN_pin_7 & CLB_2_1_IN_pin_6 & CLB_2_1_IN_pin_5 & CLB_2_1_IN_pin_4 & CLB_2_1_IN_pin_3 & CLB_2_1_IN_pin_2 & CLB_2_1_IN_pin_1 & CLB_2_1_IN_pin_0;
	CLB_2_2_inputs <= CLB_2_2_IN_pin_9 & CLB_2_2_IN_pin_8 & CLB_2_2_IN_pin_7 & CLB_2_2_IN_pin_6 & CLB_2_2_IN_pin_5 & CLB_2_2_IN_pin_4 & CLB_2_2_IN_pin_3 & CLB_2_2_IN_pin_2 & CLB_2_2_IN_pin_1 & CLB_2_2_IN_pin_0;
	CLB_2_3_inputs <= CLB_2_3_IN_pin_9 & CLB_2_3_IN_pin_8 & CLB_2_3_IN_pin_7 & CLB_2_3_IN_pin_6 & CLB_2_3_IN_pin_5 & CLB_2_3_IN_pin_4 & CLB_2_3_IN_pin_3 & CLB_2_3_IN_pin_2 & CLB_2_3_IN_pin_1 & CLB_2_3_IN_pin_0;
	CLB_2_4_inputs <= CLB_2_4_IN_pin_9 & CLB_2_4_IN_pin_8 & CLB_2_4_IN_pin_7 & CLB_2_4_IN_pin_6 & CLB_2_4_IN_pin_5 & CLB_2_4_IN_pin_4 & CLB_2_4_IN_pin_3 & CLB_2_4_IN_pin_2 & CLB_2_4_IN_pin_1 & CLB_2_4_IN_pin_0;
	CLB_2_5_inputs <= CLB_2_5_IN_pin_9 & CLB_2_5_IN_pin_8 & CLB_2_5_IN_pin_7 & CLB_2_5_IN_pin_6 & CLB_2_5_IN_pin_5 & CLB_2_5_IN_pin_4 & CLB_2_5_IN_pin_3 & CLB_2_5_IN_pin_2 & CLB_2_5_IN_pin_1 & CLB_2_5_IN_pin_0;
	CLB_2_6_inputs <= CLB_2_6_IN_pin_9 & CLB_2_6_IN_pin_8 & CLB_2_6_IN_pin_7 & CLB_2_6_IN_pin_6 & CLB_2_6_IN_pin_5 & CLB_2_6_IN_pin_4 & CLB_2_6_IN_pin_3 & CLB_2_6_IN_pin_2 & CLB_2_6_IN_pin_1 & CLB_2_6_IN_pin_0;
	CLB_3_1_inputs <= CLB_3_1_IN_pin_9 & CLB_3_1_IN_pin_8 & CLB_3_1_IN_pin_7 & CLB_3_1_IN_pin_6 & CLB_3_1_IN_pin_5 & CLB_3_1_IN_pin_4 & CLB_3_1_IN_pin_3 & CLB_3_1_IN_pin_2 & CLB_3_1_IN_pin_1 & CLB_3_1_IN_pin_0;
	CLB_3_2_inputs <= CLB_3_2_IN_pin_9 & CLB_3_2_IN_pin_8 & CLB_3_2_IN_pin_7 & CLB_3_2_IN_pin_6 & CLB_3_2_IN_pin_5 & CLB_3_2_IN_pin_4 & CLB_3_2_IN_pin_3 & CLB_3_2_IN_pin_2 & CLB_3_2_IN_pin_1 & CLB_3_2_IN_pin_0;
	CLB_3_3_inputs <= CLB_3_3_IN_pin_9 & CLB_3_3_IN_pin_8 & CLB_3_3_IN_pin_7 & CLB_3_3_IN_pin_6 & CLB_3_3_IN_pin_5 & CLB_3_3_IN_pin_4 & CLB_3_3_IN_pin_3 & CLB_3_3_IN_pin_2 & CLB_3_3_IN_pin_1 & CLB_3_3_IN_pin_0;
	CLB_3_4_inputs <= CLB_3_4_IN_pin_9 & CLB_3_4_IN_pin_8 & CLB_3_4_IN_pin_7 & CLB_3_4_IN_pin_6 & CLB_3_4_IN_pin_5 & CLB_3_4_IN_pin_4 & CLB_3_4_IN_pin_3 & CLB_3_4_IN_pin_2 & CLB_3_4_IN_pin_1 & CLB_3_4_IN_pin_0;
	CLB_3_5_inputs <= CLB_3_5_IN_pin_9 & CLB_3_5_IN_pin_8 & CLB_3_5_IN_pin_7 & CLB_3_5_IN_pin_6 & CLB_3_5_IN_pin_5 & CLB_3_5_IN_pin_4 & CLB_3_5_IN_pin_3 & CLB_3_5_IN_pin_2 & CLB_3_5_IN_pin_1 & CLB_3_5_IN_pin_0;
	CLB_3_6_inputs <= CLB_3_6_IN_pin_9 & CLB_3_6_IN_pin_8 & CLB_3_6_IN_pin_7 & CLB_3_6_IN_pin_6 & CLB_3_6_IN_pin_5 & CLB_3_6_IN_pin_4 & CLB_3_6_IN_pin_3 & CLB_3_6_IN_pin_2 & CLB_3_6_IN_pin_1 & CLB_3_6_IN_pin_0;
	CLB_4_1_inputs <= CLB_4_1_IN_pin_9 & CLB_4_1_IN_pin_8 & CLB_4_1_IN_pin_7 & CLB_4_1_IN_pin_6 & CLB_4_1_IN_pin_5 & CLB_4_1_IN_pin_4 & CLB_4_1_IN_pin_3 & CLB_4_1_IN_pin_2 & CLB_4_1_IN_pin_1 & CLB_4_1_IN_pin_0;
	CLB_4_2_inputs <= CLB_4_2_IN_pin_9 & CLB_4_2_IN_pin_8 & CLB_4_2_IN_pin_7 & CLB_4_2_IN_pin_6 & CLB_4_2_IN_pin_5 & CLB_4_2_IN_pin_4 & CLB_4_2_IN_pin_3 & CLB_4_2_IN_pin_2 & CLB_4_2_IN_pin_1 & CLB_4_2_IN_pin_0;
	CLB_4_3_inputs <= CLB_4_3_IN_pin_9 & CLB_4_3_IN_pin_8 & CLB_4_3_IN_pin_7 & CLB_4_3_IN_pin_6 & CLB_4_3_IN_pin_5 & CLB_4_3_IN_pin_4 & CLB_4_3_IN_pin_3 & CLB_4_3_IN_pin_2 & CLB_4_3_IN_pin_1 & CLB_4_3_IN_pin_0;
	CLB_4_4_inputs <= CLB_4_4_IN_pin_9 & CLB_4_4_IN_pin_8 & CLB_4_4_IN_pin_7 & CLB_4_4_IN_pin_6 & CLB_4_4_IN_pin_5 & CLB_4_4_IN_pin_4 & CLB_4_4_IN_pin_3 & CLB_4_4_IN_pin_2 & CLB_4_4_IN_pin_1 & CLB_4_4_IN_pin_0;
	CLB_4_5_inputs <= CLB_4_5_IN_pin_9 & CLB_4_5_IN_pin_8 & CLB_4_5_IN_pin_7 & CLB_4_5_IN_pin_6 & CLB_4_5_IN_pin_5 & CLB_4_5_IN_pin_4 & CLB_4_5_IN_pin_3 & CLB_4_5_IN_pin_2 & CLB_4_5_IN_pin_1 & CLB_4_5_IN_pin_0;
	CLB_4_6_inputs <= CLB_4_6_IN_pin_9 & CLB_4_6_IN_pin_8 & CLB_4_6_IN_pin_7 & CLB_4_6_IN_pin_6 & CLB_4_6_IN_pin_5 & CLB_4_6_IN_pin_4 & CLB_4_6_IN_pin_3 & CLB_4_6_IN_pin_2 & CLB_4_6_IN_pin_1 & CLB_4_6_IN_pin_0;
	CLB_5_1_inputs <= CLB_5_1_IN_pin_9 & CLB_5_1_IN_pin_8 & CLB_5_1_IN_pin_7 & CLB_5_1_IN_pin_6 & CLB_5_1_IN_pin_5 & CLB_5_1_IN_pin_4 & CLB_5_1_IN_pin_3 & CLB_5_1_IN_pin_2 & CLB_5_1_IN_pin_1 & CLB_5_1_IN_pin_0;
	CLB_5_2_inputs <= CLB_5_2_IN_pin_9 & CLB_5_2_IN_pin_8 & CLB_5_2_IN_pin_7 & CLB_5_2_IN_pin_6 & CLB_5_2_IN_pin_5 & CLB_5_2_IN_pin_4 & CLB_5_2_IN_pin_3 & CLB_5_2_IN_pin_2 & CLB_5_2_IN_pin_1 & CLB_5_2_IN_pin_0;
	CLB_5_3_inputs <= CLB_5_3_IN_pin_9 & CLB_5_3_IN_pin_8 & CLB_5_3_IN_pin_7 & CLB_5_3_IN_pin_6 & CLB_5_3_IN_pin_5 & CLB_5_3_IN_pin_4 & CLB_5_3_IN_pin_3 & CLB_5_3_IN_pin_2 & CLB_5_3_IN_pin_1 & CLB_5_3_IN_pin_0;
	CLB_5_4_inputs <= CLB_5_4_IN_pin_9 & CLB_5_4_IN_pin_8 & CLB_5_4_IN_pin_7 & CLB_5_4_IN_pin_6 & CLB_5_4_IN_pin_5 & CLB_5_4_IN_pin_4 & CLB_5_4_IN_pin_3 & CLB_5_4_IN_pin_2 & CLB_5_4_IN_pin_1 & CLB_5_4_IN_pin_0;
	CLB_5_5_inputs <= CLB_5_5_IN_pin_9 & CLB_5_5_IN_pin_8 & CLB_5_5_IN_pin_7 & CLB_5_5_IN_pin_6 & CLB_5_5_IN_pin_5 & CLB_5_5_IN_pin_4 & CLB_5_5_IN_pin_3 & CLB_5_5_IN_pin_2 & CLB_5_5_IN_pin_1 & CLB_5_5_IN_pin_0;
	CLB_5_6_inputs <= CLB_5_6_IN_pin_9 & CLB_5_6_IN_pin_8 & CLB_5_6_IN_pin_7 & CLB_5_6_IN_pin_6 & CLB_5_6_IN_pin_5 & CLB_5_6_IN_pin_4 & CLB_5_6_IN_pin_3 & CLB_5_6_IN_pin_2 & CLB_5_6_IN_pin_1 & CLB_5_6_IN_pin_0;
	CLB_6_1_inputs <= CLB_6_1_IN_pin_9 & CLB_6_1_IN_pin_8 & CLB_6_1_IN_pin_7 & CLB_6_1_IN_pin_6 & CLB_6_1_IN_pin_5 & CLB_6_1_IN_pin_4 & CLB_6_1_IN_pin_3 & CLB_6_1_IN_pin_2 & CLB_6_1_IN_pin_1 & CLB_6_1_IN_pin_0;
	CLB_6_2_inputs <= CLB_6_2_IN_pin_9 & CLB_6_2_IN_pin_8 & CLB_6_2_IN_pin_7 & CLB_6_2_IN_pin_6 & CLB_6_2_IN_pin_5 & CLB_6_2_IN_pin_4 & CLB_6_2_IN_pin_3 & CLB_6_2_IN_pin_2 & CLB_6_2_IN_pin_1 & CLB_6_2_IN_pin_0;
	CLB_6_3_inputs <= CLB_6_3_IN_pin_9 & CLB_6_3_IN_pin_8 & CLB_6_3_IN_pin_7 & CLB_6_3_IN_pin_6 & CLB_6_3_IN_pin_5 & CLB_6_3_IN_pin_4 & CLB_6_3_IN_pin_3 & CLB_6_3_IN_pin_2 & CLB_6_3_IN_pin_1 & CLB_6_3_IN_pin_0;
	CLB_6_4_inputs <= CLB_6_4_IN_pin_9 & CLB_6_4_IN_pin_8 & CLB_6_4_IN_pin_7 & CLB_6_4_IN_pin_6 & CLB_6_4_IN_pin_5 & CLB_6_4_IN_pin_4 & CLB_6_4_IN_pin_3 & CLB_6_4_IN_pin_2 & CLB_6_4_IN_pin_1 & CLB_6_4_IN_pin_0;
	CLB_6_5_inputs <= CLB_6_5_IN_pin_9 & CLB_6_5_IN_pin_8 & CLB_6_5_IN_pin_7 & CLB_6_5_IN_pin_6 & CLB_6_5_IN_pin_5 & CLB_6_5_IN_pin_4 & CLB_6_5_IN_pin_3 & CLB_6_5_IN_pin_2 & CLB_6_5_IN_pin_1 & CLB_6_5_IN_pin_0;
	CLB_6_6_inputs <= CLB_6_6_IN_pin_9 & CLB_6_6_IN_pin_8 & CLB_6_6_IN_pin_7 & CLB_6_6_IN_pin_6 & CLB_6_6_IN_pin_5 & CLB_6_6_IN_pin_4 & CLB_6_6_IN_pin_3 & CLB_6_6_IN_pin_2 & CLB_6_6_IN_pin_1 & CLB_6_6_IN_pin_0;
	CLB_7_1_inputs <= CLB_7_1_IN_pin_9 & CLB_7_1_IN_pin_8 & CLB_7_1_IN_pin_7 & CLB_7_1_IN_pin_6 & CLB_7_1_IN_pin_5 & CLB_7_1_IN_pin_4 & CLB_7_1_IN_pin_3 & CLB_7_1_IN_pin_2 & CLB_7_1_IN_pin_1 & CLB_7_1_IN_pin_0;
	CLB_7_2_inputs <= CLB_7_2_IN_pin_9 & CLB_7_2_IN_pin_8 & CLB_7_2_IN_pin_7 & CLB_7_2_IN_pin_6 & CLB_7_2_IN_pin_5 & CLB_7_2_IN_pin_4 & CLB_7_2_IN_pin_3 & CLB_7_2_IN_pin_2 & CLB_7_2_IN_pin_1 & CLB_7_2_IN_pin_0;
	CLB_7_3_inputs <= CLB_7_3_IN_pin_9 & CLB_7_3_IN_pin_8 & CLB_7_3_IN_pin_7 & CLB_7_3_IN_pin_6 & CLB_7_3_IN_pin_5 & CLB_7_3_IN_pin_4 & CLB_7_3_IN_pin_3 & CLB_7_3_IN_pin_2 & CLB_7_3_IN_pin_1 & CLB_7_3_IN_pin_0;
	CLB_7_4_inputs <= CLB_7_4_IN_pin_9 & CLB_7_4_IN_pin_8 & CLB_7_4_IN_pin_7 & CLB_7_4_IN_pin_6 & CLB_7_4_IN_pin_5 & CLB_7_4_IN_pin_4 & CLB_7_4_IN_pin_3 & CLB_7_4_IN_pin_2 & CLB_7_4_IN_pin_1 & CLB_7_4_IN_pin_0;
	CLB_7_5_inputs <= CLB_7_5_IN_pin_9 & CLB_7_5_IN_pin_8 & CLB_7_5_IN_pin_7 & CLB_7_5_IN_pin_6 & CLB_7_5_IN_pin_5 & CLB_7_5_IN_pin_4 & CLB_7_5_IN_pin_3 & CLB_7_5_IN_pin_2 & CLB_7_5_IN_pin_1 & CLB_7_5_IN_pin_0;
	CLB_7_6_inputs <= CLB_7_6_IN_pin_9 & CLB_7_6_IN_pin_8 & CLB_7_6_IN_pin_7 & CLB_7_6_IN_pin_6 & CLB_7_6_IN_pin_5 & CLB_7_6_IN_pin_4 & CLB_7_6_IN_pin_3 & CLB_7_6_IN_pin_2 & CLB_7_6_IN_pin_1 & CLB_7_6_IN_pin_0;
	CLB_8_1_inputs <= CLB_8_1_IN_pin_9 & CLB_8_1_IN_pin_8 & CLB_8_1_IN_pin_7 & CLB_8_1_IN_pin_6 & CLB_8_1_IN_pin_5 & CLB_8_1_IN_pin_4 & CLB_8_1_IN_pin_3 & CLB_8_1_IN_pin_2 & CLB_8_1_IN_pin_1 & CLB_8_1_IN_pin_0;
	CLB_8_2_inputs <= CLB_8_2_IN_pin_9 & CLB_8_2_IN_pin_8 & CLB_8_2_IN_pin_7 & CLB_8_2_IN_pin_6 & CLB_8_2_IN_pin_5 & CLB_8_2_IN_pin_4 & CLB_8_2_IN_pin_3 & CLB_8_2_IN_pin_2 & CLB_8_2_IN_pin_1 & CLB_8_2_IN_pin_0;
	CLB_8_3_inputs <= CLB_8_3_IN_pin_9 & CLB_8_3_IN_pin_8 & CLB_8_3_IN_pin_7 & CLB_8_3_IN_pin_6 & CLB_8_3_IN_pin_5 & CLB_8_3_IN_pin_4 & CLB_8_3_IN_pin_3 & CLB_8_3_IN_pin_2 & CLB_8_3_IN_pin_1 & CLB_8_3_IN_pin_0;
	CLB_8_4_inputs <= CLB_8_4_IN_pin_9 & CLB_8_4_IN_pin_8 & CLB_8_4_IN_pin_7 & CLB_8_4_IN_pin_6 & CLB_8_4_IN_pin_5 & CLB_8_4_IN_pin_4 & CLB_8_4_IN_pin_3 & CLB_8_4_IN_pin_2 & CLB_8_4_IN_pin_1 & CLB_8_4_IN_pin_0;
	CLB_8_5_inputs <= CLB_8_5_IN_pin_9 & CLB_8_5_IN_pin_8 & CLB_8_5_IN_pin_7 & CLB_8_5_IN_pin_6 & CLB_8_5_IN_pin_5 & CLB_8_5_IN_pin_4 & CLB_8_5_IN_pin_3 & CLB_8_5_IN_pin_2 & CLB_8_5_IN_pin_1 & CLB_8_5_IN_pin_0;
	CLB_8_6_inputs <= CLB_8_6_IN_pin_9 & CLB_8_6_IN_pin_8 & CLB_8_6_IN_pin_7 & CLB_8_6_IN_pin_6 & CLB_8_6_IN_pin_5 & CLB_8_6_IN_pin_4 & CLB_8_6_IN_pin_3 & CLB_8_6_IN_pin_2 & CLB_8_6_IN_pin_1 & CLB_8_6_IN_pin_0;

	-- CLB outputs --
	CLB_1_1_OUT_pin_0 <= CLB_1_1_outputs(0);
	CLB_1_1_OUT_pin_1 <= CLB_1_1_outputs(1);
	CLB_1_1_OUT_pin_2 <= CLB_1_1_outputs(2);
	CLB_1_1_OUT_pin_3 <= CLB_1_1_outputs(3);
	CLB_1_2_OUT_pin_0 <= CLB_1_2_outputs(0);
	CLB_1_2_OUT_pin_1 <= CLB_1_2_outputs(1);
	CLB_1_2_OUT_pin_2 <= CLB_1_2_outputs(2);
	CLB_1_2_OUT_pin_3 <= CLB_1_2_outputs(3);
	CLB_1_3_OUT_pin_0 <= CLB_1_3_outputs(0);
	CLB_1_3_OUT_pin_1 <= CLB_1_3_outputs(1);
	CLB_1_3_OUT_pin_2 <= CLB_1_3_outputs(2);
	CLB_1_3_OUT_pin_3 <= CLB_1_3_outputs(3);
	CLB_1_4_OUT_pin_0 <= CLB_1_4_outputs(0);
	CLB_1_4_OUT_pin_1 <= CLB_1_4_outputs(1);
	CLB_1_4_OUT_pin_2 <= CLB_1_4_outputs(2);
	CLB_1_4_OUT_pin_3 <= CLB_1_4_outputs(3);
	CLB_1_5_OUT_pin_0 <= CLB_1_5_outputs(0);
	CLB_1_5_OUT_pin_1 <= CLB_1_5_outputs(1);
	CLB_1_5_OUT_pin_2 <= CLB_1_5_outputs(2);
	CLB_1_5_OUT_pin_3 <= CLB_1_5_outputs(3);
	CLB_1_6_OUT_pin_0 <= CLB_1_6_outputs(0);
	CLB_1_6_OUT_pin_1 <= CLB_1_6_outputs(1);
	CLB_1_6_OUT_pin_2 <= CLB_1_6_outputs(2);
	CLB_1_6_OUT_pin_3 <= CLB_1_6_outputs(3);
	CLB_2_1_OUT_pin_0 <= CLB_2_1_outputs(0);
	CLB_2_1_OUT_pin_1 <= CLB_2_1_outputs(1);
	CLB_2_1_OUT_pin_2 <= CLB_2_1_outputs(2);
	CLB_2_1_OUT_pin_3 <= CLB_2_1_outputs(3);
	CLB_2_2_OUT_pin_0 <= CLB_2_2_outputs(0);
	CLB_2_2_OUT_pin_1 <= CLB_2_2_outputs(1);
	CLB_2_2_OUT_pin_2 <= CLB_2_2_outputs(2);
	CLB_2_2_OUT_pin_3 <= CLB_2_2_outputs(3);
	CLB_2_3_OUT_pin_0 <= CLB_2_3_outputs(0);
	CLB_2_3_OUT_pin_1 <= CLB_2_3_outputs(1);
	CLB_2_3_OUT_pin_2 <= CLB_2_3_outputs(2);
	CLB_2_3_OUT_pin_3 <= CLB_2_3_outputs(3);
	CLB_2_4_OUT_pin_0 <= CLB_2_4_outputs(0);
	CLB_2_4_OUT_pin_1 <= CLB_2_4_outputs(1);
	CLB_2_4_OUT_pin_2 <= CLB_2_4_outputs(2);
	CLB_2_4_OUT_pin_3 <= CLB_2_4_outputs(3);
	CLB_2_5_OUT_pin_0 <= CLB_2_5_outputs(0);
	CLB_2_5_OUT_pin_1 <= CLB_2_5_outputs(1);
	CLB_2_5_OUT_pin_2 <= CLB_2_5_outputs(2);
	CLB_2_5_OUT_pin_3 <= CLB_2_5_outputs(3);
	CLB_2_6_OUT_pin_0 <= CLB_2_6_outputs(0);
	CLB_2_6_OUT_pin_1 <= CLB_2_6_outputs(1);
	CLB_2_6_OUT_pin_2 <= CLB_2_6_outputs(2);
	CLB_2_6_OUT_pin_3 <= CLB_2_6_outputs(3);
	CLB_3_1_OUT_pin_0 <= CLB_3_1_outputs(0);
	CLB_3_1_OUT_pin_1 <= CLB_3_1_outputs(1);
	CLB_3_1_OUT_pin_2 <= CLB_3_1_outputs(2);
	CLB_3_1_OUT_pin_3 <= CLB_3_1_outputs(3);
	CLB_3_2_OUT_pin_0 <= CLB_3_2_outputs(0);
	CLB_3_2_OUT_pin_1 <= CLB_3_2_outputs(1);
	CLB_3_2_OUT_pin_2 <= CLB_3_2_outputs(2);
	CLB_3_2_OUT_pin_3 <= CLB_3_2_outputs(3);
	CLB_3_3_OUT_pin_0 <= CLB_3_3_outputs(0);
	CLB_3_3_OUT_pin_1 <= CLB_3_3_outputs(1);
	CLB_3_3_OUT_pin_2 <= CLB_3_3_outputs(2);
	CLB_3_3_OUT_pin_3 <= CLB_3_3_outputs(3);
	CLB_3_4_OUT_pin_0 <= CLB_3_4_outputs(0);
	CLB_3_4_OUT_pin_1 <= CLB_3_4_outputs(1);
	CLB_3_4_OUT_pin_2 <= CLB_3_4_outputs(2);
	CLB_3_4_OUT_pin_3 <= CLB_3_4_outputs(3);
	CLB_3_5_OUT_pin_0 <= CLB_3_5_outputs(0);
	CLB_3_5_OUT_pin_1 <= CLB_3_5_outputs(1);
	CLB_3_5_OUT_pin_2 <= CLB_3_5_outputs(2);
	CLB_3_5_OUT_pin_3 <= CLB_3_5_outputs(3);
	CLB_3_6_OUT_pin_0 <= CLB_3_6_outputs(0);
	CLB_3_6_OUT_pin_1 <= CLB_3_6_outputs(1);
	CLB_3_6_OUT_pin_2 <= CLB_3_6_outputs(2);
	CLB_3_6_OUT_pin_3 <= CLB_3_6_outputs(3);
	CLB_4_1_OUT_pin_0 <= CLB_4_1_outputs(0);
	CLB_4_1_OUT_pin_1 <= CLB_4_1_outputs(1);
	CLB_4_1_OUT_pin_2 <= CLB_4_1_outputs(2);
	CLB_4_1_OUT_pin_3 <= CLB_4_1_outputs(3);
	CLB_4_2_OUT_pin_0 <= CLB_4_2_outputs(0);
	CLB_4_2_OUT_pin_1 <= CLB_4_2_outputs(1);
	CLB_4_2_OUT_pin_2 <= CLB_4_2_outputs(2);
	CLB_4_2_OUT_pin_3 <= CLB_4_2_outputs(3);
	CLB_4_3_OUT_pin_0 <= CLB_4_3_outputs(0);
	CLB_4_3_OUT_pin_1 <= CLB_4_3_outputs(1);
	CLB_4_3_OUT_pin_2 <= CLB_4_3_outputs(2);
	CLB_4_3_OUT_pin_3 <= CLB_4_3_outputs(3);
	CLB_4_4_OUT_pin_0 <= CLB_4_4_outputs(0);
	CLB_4_4_OUT_pin_1 <= CLB_4_4_outputs(1);
	CLB_4_4_OUT_pin_2 <= CLB_4_4_outputs(2);
	CLB_4_4_OUT_pin_3 <= CLB_4_4_outputs(3);
	CLB_4_5_OUT_pin_0 <= CLB_4_5_outputs(0);
	CLB_4_5_OUT_pin_1 <= CLB_4_5_outputs(1);
	CLB_4_5_OUT_pin_2 <= CLB_4_5_outputs(2);
	CLB_4_5_OUT_pin_3 <= CLB_4_5_outputs(3);
	CLB_4_6_OUT_pin_0 <= CLB_4_6_outputs(0);
	CLB_4_6_OUT_pin_1 <= CLB_4_6_outputs(1);
	CLB_4_6_OUT_pin_2 <= CLB_4_6_outputs(2);
	CLB_4_6_OUT_pin_3 <= CLB_4_6_outputs(3);
	CLB_5_1_OUT_pin_0 <= CLB_5_1_outputs(0);
	CLB_5_1_OUT_pin_1 <= CLB_5_1_outputs(1);
	CLB_5_1_OUT_pin_2 <= CLB_5_1_outputs(2);
	CLB_5_1_OUT_pin_3 <= CLB_5_1_outputs(3);
	CLB_5_2_OUT_pin_0 <= CLB_5_2_outputs(0);
	CLB_5_2_OUT_pin_1 <= CLB_5_2_outputs(1);
	CLB_5_2_OUT_pin_2 <= CLB_5_2_outputs(2);
	CLB_5_2_OUT_pin_3 <= CLB_5_2_outputs(3);
	CLB_5_3_OUT_pin_0 <= CLB_5_3_outputs(0);
	CLB_5_3_OUT_pin_1 <= CLB_5_3_outputs(1);
	CLB_5_3_OUT_pin_2 <= CLB_5_3_outputs(2);
	CLB_5_3_OUT_pin_3 <= CLB_5_3_outputs(3);
	CLB_5_4_OUT_pin_0 <= CLB_5_4_outputs(0);
	CLB_5_4_OUT_pin_1 <= CLB_5_4_outputs(1);
	CLB_5_4_OUT_pin_2 <= CLB_5_4_outputs(2);
	CLB_5_4_OUT_pin_3 <= CLB_5_4_outputs(3);
	CLB_5_5_OUT_pin_0 <= CLB_5_5_outputs(0);
	CLB_5_5_OUT_pin_1 <= CLB_5_5_outputs(1);
	CLB_5_5_OUT_pin_2 <= CLB_5_5_outputs(2);
	CLB_5_5_OUT_pin_3 <= CLB_5_5_outputs(3);
	CLB_5_6_OUT_pin_0 <= CLB_5_6_outputs(0);
	CLB_5_6_OUT_pin_1 <= CLB_5_6_outputs(1);
	CLB_5_6_OUT_pin_2 <= CLB_5_6_outputs(2);
	CLB_5_6_OUT_pin_3 <= CLB_5_6_outputs(3);
	CLB_6_1_OUT_pin_0 <= CLB_6_1_outputs(0);
	CLB_6_1_OUT_pin_1 <= CLB_6_1_outputs(1);
	CLB_6_1_OUT_pin_2 <= CLB_6_1_outputs(2);
	CLB_6_1_OUT_pin_3 <= CLB_6_1_outputs(3);
	CLB_6_2_OUT_pin_0 <= CLB_6_2_outputs(0);
	CLB_6_2_OUT_pin_1 <= CLB_6_2_outputs(1);
	CLB_6_2_OUT_pin_2 <= CLB_6_2_outputs(2);
	CLB_6_2_OUT_pin_3 <= CLB_6_2_outputs(3);
	CLB_6_3_OUT_pin_0 <= CLB_6_3_outputs(0);
	CLB_6_3_OUT_pin_1 <= CLB_6_3_outputs(1);
	CLB_6_3_OUT_pin_2 <= CLB_6_3_outputs(2);
	CLB_6_3_OUT_pin_3 <= CLB_6_3_outputs(3);
	CLB_6_4_OUT_pin_0 <= CLB_6_4_outputs(0);
	CLB_6_4_OUT_pin_1 <= CLB_6_4_outputs(1);
	CLB_6_4_OUT_pin_2 <= CLB_6_4_outputs(2);
	CLB_6_4_OUT_pin_3 <= CLB_6_4_outputs(3);
	CLB_6_5_OUT_pin_0 <= CLB_6_5_outputs(0);
	CLB_6_5_OUT_pin_1 <= CLB_6_5_outputs(1);
	CLB_6_5_OUT_pin_2 <= CLB_6_5_outputs(2);
	CLB_6_5_OUT_pin_3 <= CLB_6_5_outputs(3);
	CLB_6_6_OUT_pin_0 <= CLB_6_6_outputs(0);
	CLB_6_6_OUT_pin_1 <= CLB_6_6_outputs(1);
	CLB_6_6_OUT_pin_2 <= CLB_6_6_outputs(2);
	CLB_6_6_OUT_pin_3 <= CLB_6_6_outputs(3);
	CLB_7_1_OUT_pin_0 <= CLB_7_1_outputs(0);
	CLB_7_1_OUT_pin_1 <= CLB_7_1_outputs(1);
	CLB_7_1_OUT_pin_2 <= CLB_7_1_outputs(2);
	CLB_7_1_OUT_pin_3 <= CLB_7_1_outputs(3);
	CLB_7_2_OUT_pin_0 <= CLB_7_2_outputs(0);
	CLB_7_2_OUT_pin_1 <= CLB_7_2_outputs(1);
	CLB_7_2_OUT_pin_2 <= CLB_7_2_outputs(2);
	CLB_7_2_OUT_pin_3 <= CLB_7_2_outputs(3);
	CLB_7_3_OUT_pin_0 <= CLB_7_3_outputs(0);
	CLB_7_3_OUT_pin_1 <= CLB_7_3_outputs(1);
	CLB_7_3_OUT_pin_2 <= CLB_7_3_outputs(2);
	CLB_7_3_OUT_pin_3 <= CLB_7_3_outputs(3);
	CLB_7_4_OUT_pin_0 <= CLB_7_4_outputs(0);
	CLB_7_4_OUT_pin_1 <= CLB_7_4_outputs(1);
	CLB_7_4_OUT_pin_2 <= CLB_7_4_outputs(2);
	CLB_7_4_OUT_pin_3 <= CLB_7_4_outputs(3);
	CLB_7_5_OUT_pin_0 <= CLB_7_5_outputs(0);
	CLB_7_5_OUT_pin_1 <= CLB_7_5_outputs(1);
	CLB_7_5_OUT_pin_2 <= CLB_7_5_outputs(2);
	CLB_7_5_OUT_pin_3 <= CLB_7_5_outputs(3);
	CLB_7_6_OUT_pin_0 <= CLB_7_6_outputs(0);
	CLB_7_6_OUT_pin_1 <= CLB_7_6_outputs(1);
	CLB_7_6_OUT_pin_2 <= CLB_7_6_outputs(2);
	CLB_7_6_OUT_pin_3 <= CLB_7_6_outputs(3);
	CLB_8_1_OUT_pin_0 <= CLB_8_1_outputs(0);
	CLB_8_1_OUT_pin_1 <= CLB_8_1_outputs(1);
	CLB_8_1_OUT_pin_2 <= CLB_8_1_outputs(2);
	CLB_8_1_OUT_pin_3 <= CLB_8_1_outputs(3);
	CLB_8_2_OUT_pin_0 <= CLB_8_2_outputs(0);
	CLB_8_2_OUT_pin_1 <= CLB_8_2_outputs(1);
	CLB_8_2_OUT_pin_2 <= CLB_8_2_outputs(2);
	CLB_8_2_OUT_pin_3 <= CLB_8_2_outputs(3);
	CLB_8_3_OUT_pin_0 <= CLB_8_3_outputs(0);
	CLB_8_3_OUT_pin_1 <= CLB_8_3_outputs(1);
	CLB_8_3_OUT_pin_2 <= CLB_8_3_outputs(2);
	CLB_8_3_OUT_pin_3 <= CLB_8_3_outputs(3);
	CLB_8_4_OUT_pin_0 <= CLB_8_4_outputs(0);
	CLB_8_4_OUT_pin_1 <= CLB_8_4_outputs(1);
	CLB_8_4_OUT_pin_2 <= CLB_8_4_outputs(2);
	CLB_8_4_OUT_pin_3 <= CLB_8_4_outputs(3);
	CLB_8_5_OUT_pin_0 <= CLB_8_5_outputs(0);
	CLB_8_5_OUT_pin_1 <= CLB_8_5_outputs(1);
	CLB_8_5_OUT_pin_2 <= CLB_8_5_outputs(2);
	CLB_8_5_OUT_pin_3 <= CLB_8_5_outputs(3);
	CLB_8_6_OUT_pin_0 <= CLB_8_6_outputs(0);
	CLB_8_6_OUT_pin_1 <= CLB_8_6_outputs(1);
	CLB_8_6_OUT_pin_2 <= CLB_8_6_outputs(2);
	CLB_8_6_OUT_pin_3 <= CLB_8_6_outputs(3);

	-- CLB snapshot out --
	snap_out(  3 downto   0) <= CLB_1_1_snapshot_out;
	snap_out(  7 downto   4) <= CLB_1_2_snapshot_out;
	snap_out( 11 downto   8) <= CLB_1_3_snapshot_out;
	snap_out( 15 downto  12) <= CLB_1_4_snapshot_out;
	snap_out( 19 downto  16) <= CLB_1_5_snapshot_out;
	snap_out( 23 downto  20) <= CLB_1_6_snapshot_out;
	snap_out( 27 downto  24) <= CLB_2_1_snapshot_out;
	snap_out( 31 downto  28) <= CLB_2_2_snapshot_out;
	snap_out( 35 downto  32) <= CLB_2_3_snapshot_out;
	snap_out( 39 downto  36) <= CLB_2_4_snapshot_out;
	snap_out( 43 downto  40) <= CLB_2_5_snapshot_out;
	snap_out( 47 downto  44) <= CLB_2_6_snapshot_out;
	snap_out( 51 downto  48) <= CLB_3_1_snapshot_out;
	snap_out( 55 downto  52) <= CLB_3_2_snapshot_out;
	snap_out( 59 downto  56) <= CLB_3_3_snapshot_out;
	snap_out( 63 downto  60) <= CLB_3_4_snapshot_out;
	snap_out( 67 downto  64) <= CLB_3_5_snapshot_out;
	snap_out( 71 downto  68) <= CLB_3_6_snapshot_out;
	snap_out( 75 downto  72) <= CLB_4_1_snapshot_out;
	snap_out( 79 downto  76) <= CLB_4_2_snapshot_out;
	snap_out( 83 downto  80) <= CLB_4_3_snapshot_out;
	snap_out( 87 downto  84) <= CLB_4_4_snapshot_out;
	snap_out( 91 downto  88) <= CLB_4_5_snapshot_out;
	snap_out( 95 downto  92) <= CLB_4_6_snapshot_out;
	snap_out( 99 downto  96) <= CLB_5_1_snapshot_out;
	snap_out(103 downto 100) <= CLB_5_2_snapshot_out;
	snap_out(107 downto 104) <= CLB_5_3_snapshot_out;
	snap_out(111 downto 108) <= CLB_5_4_snapshot_out;
	snap_out(115 downto 112) <= CLB_5_5_snapshot_out;
	snap_out(119 downto 116) <= CLB_5_6_snapshot_out;
	snap_out(123 downto 120) <= CLB_6_1_snapshot_out;
	snap_out(127 downto 124) <= CLB_6_2_snapshot_out;
	snap_out(131 downto 128) <= CLB_6_3_snapshot_out;
	snap_out(135 downto 132) <= CLB_6_4_snapshot_out;
	snap_out(139 downto 136) <= CLB_6_5_snapshot_out;
	snap_out(143 downto 140) <= CLB_6_6_snapshot_out;
	snap_out(147 downto 144) <= CLB_7_1_snapshot_out;
	snap_out(151 downto 148) <= CLB_7_2_snapshot_out;
	snap_out(155 downto 152) <= CLB_7_3_snapshot_out;
	snap_out(159 downto 156) <= CLB_7_4_snapshot_out;
	snap_out(163 downto 160) <= CLB_7_5_snapshot_out;
	snap_out(167 downto 164) <= CLB_7_6_snapshot_out;
	snap_out(171 downto 168) <= CLB_8_1_snapshot_out;
	snap_out(175 downto 172) <= CLB_8_2_snapshot_out;
	snap_out(179 downto 176) <= CLB_8_3_snapshot_out;
	snap_out(183 downto 180) <= CLB_8_4_snapshot_out;
	snap_out(187 downto 184) <= CLB_8_5_snapshot_out;
	snap_out(191 downto 188) <= CLB_8_6_snapshot_out;

	-- CLB instanciations --

	CLB_1_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(3 downto 0),
	           snap_out     => CLB_1_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(131 downto 0),
	           inputs       => CLB_1_1_inputs,
	           outputs      => CLB_1_1_outputs);
	
	CLB_1_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(7 downto 4),
	           snap_out     => CLB_1_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(263 downto 132),
	           inputs       => CLB_1_2_inputs,
	           outputs      => CLB_1_2_outputs);
	
	CLB_1_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(11 downto 8),
	           snap_out     => CLB_1_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(395 downto 264),
	           inputs       => CLB_1_3_inputs,
	           outputs      => CLB_1_3_outputs);
	
	CLB_1_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(15 downto 12),
	           snap_out     => CLB_1_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(527 downto 396),
	           inputs       => CLB_1_4_inputs,
	           outputs      => CLB_1_4_outputs);
	
	CLB_1_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(19 downto 16),
	           snap_out     => CLB_1_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(659 downto 528),
	           inputs       => CLB_1_5_inputs,
	           outputs      => CLB_1_5_outputs);
	
	CLB_1_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(23 downto 20),
	           snap_out     => CLB_1_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(791 downto 660),
	           inputs       => CLB_1_6_inputs,
	           outputs      => CLB_1_6_outputs);
	
	CLB_2_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(27 downto 24),
	           snap_out     => CLB_2_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(923 downto 792),
	           inputs       => CLB_2_1_inputs,
	           outputs      => CLB_2_1_outputs);
	
	CLB_2_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(31 downto 28),
	           snap_out     => CLB_2_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1055 downto 924),
	           inputs       => CLB_2_2_inputs,
	           outputs      => CLB_2_2_outputs);
	
	CLB_2_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(35 downto 32),
	           snap_out     => CLB_2_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1187 downto 1056),
	           inputs       => CLB_2_3_inputs,
	           outputs      => CLB_2_3_outputs);
	
	CLB_2_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(39 downto 36),
	           snap_out     => CLB_2_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1319 downto 1188),
	           inputs       => CLB_2_4_inputs,
	           outputs      => CLB_2_4_outputs);
	
	CLB_2_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(43 downto 40),
	           snap_out     => CLB_2_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1451 downto 1320),
	           inputs       => CLB_2_5_inputs,
	           outputs      => CLB_2_5_outputs);
	
	CLB_2_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(47 downto 44),
	           snap_out     => CLB_2_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1583 downto 1452),
	           inputs       => CLB_2_6_inputs,
	           outputs      => CLB_2_6_outputs);
	
	CLB_3_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(51 downto 48),
	           snap_out     => CLB_3_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1715 downto 1584),
	           inputs       => CLB_3_1_inputs,
	           outputs      => CLB_3_1_outputs);
	
	CLB_3_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(55 downto 52),
	           snap_out     => CLB_3_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1847 downto 1716),
	           inputs       => CLB_3_2_inputs,
	           outputs      => CLB_3_2_outputs);
	
	CLB_3_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(59 downto 56),
	           snap_out     => CLB_3_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(1979 downto 1848),
	           inputs       => CLB_3_3_inputs,
	           outputs      => CLB_3_3_outputs);
	
	CLB_3_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(63 downto 60),
	           snap_out     => CLB_3_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2111 downto 1980),
	           inputs       => CLB_3_4_inputs,
	           outputs      => CLB_3_4_outputs);
	
	CLB_3_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(67 downto 64),
	           snap_out     => CLB_3_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2243 downto 2112),
	           inputs       => CLB_3_5_inputs,
	           outputs      => CLB_3_5_outputs);
	
	CLB_3_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(71 downto 68),
	           snap_out     => CLB_3_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2375 downto 2244),
	           inputs       => CLB_3_6_inputs,
	           outputs      => CLB_3_6_outputs);
	
	CLB_4_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(75 downto 72),
	           snap_out     => CLB_4_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2507 downto 2376),
	           inputs       => CLB_4_1_inputs,
	           outputs      => CLB_4_1_outputs);
	
	CLB_4_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(79 downto 76),
	           snap_out     => CLB_4_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2639 downto 2508),
	           inputs       => CLB_4_2_inputs,
	           outputs      => CLB_4_2_outputs);
	
	CLB_4_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(83 downto 80),
	           snap_out     => CLB_4_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2771 downto 2640),
	           inputs       => CLB_4_3_inputs,
	           outputs      => CLB_4_3_outputs);
	
	CLB_4_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(87 downto 84),
	           snap_out     => CLB_4_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(2903 downto 2772),
	           inputs       => CLB_4_4_inputs,
	           outputs      => CLB_4_4_outputs);
	
	CLB_4_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(91 downto 88),
	           snap_out     => CLB_4_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3035 downto 2904),
	           inputs       => CLB_4_5_inputs,
	           outputs      => CLB_4_5_outputs);
	
	CLB_4_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(95 downto 92),
	           snap_out     => CLB_4_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3167 downto 3036),
	           inputs       => CLB_4_6_inputs,
	           outputs      => CLB_4_6_outputs);
	
	CLB_5_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(99 downto 96),
	           snap_out     => CLB_5_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3299 downto 3168),
	           inputs       => CLB_5_1_inputs,
	           outputs      => CLB_5_1_outputs);
	
	CLB_5_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(103 downto 100),
	           snap_out     => CLB_5_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3431 downto 3300),
	           inputs       => CLB_5_2_inputs,
	           outputs      => CLB_5_2_outputs);
	
	CLB_5_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(107 downto 104),
	           snap_out     => CLB_5_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3563 downto 3432),
	           inputs       => CLB_5_3_inputs,
	           outputs      => CLB_5_3_outputs);
	
	CLB_5_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(111 downto 108),
	           snap_out     => CLB_5_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3695 downto 3564),
	           inputs       => CLB_5_4_inputs,
	           outputs      => CLB_5_4_outputs);
	
	CLB_5_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(115 downto 112),
	           snap_out     => CLB_5_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3827 downto 3696),
	           inputs       => CLB_5_5_inputs,
	           outputs      => CLB_5_5_outputs);
	
	CLB_5_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(119 downto 116),
	           snap_out     => CLB_5_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(3959 downto 3828),
	           inputs       => CLB_5_6_inputs,
	           outputs      => CLB_5_6_outputs);
	
	CLB_6_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(123 downto 120),
	           snap_out     => CLB_6_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4091 downto 3960),
	           inputs       => CLB_6_1_inputs,
	           outputs      => CLB_6_1_outputs);
	
	CLB_6_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(127 downto 124),
	           snap_out     => CLB_6_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4223 downto 4092),
	           inputs       => CLB_6_2_inputs,
	           outputs      => CLB_6_2_outputs);
	
	CLB_6_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(131 downto 128),
	           snap_out     => CLB_6_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4355 downto 4224),
	           inputs       => CLB_6_3_inputs,
	           outputs      => CLB_6_3_outputs);
	
	CLB_6_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(135 downto 132),
	           snap_out     => CLB_6_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4487 downto 4356),
	           inputs       => CLB_6_4_inputs,
	           outputs      => CLB_6_4_outputs);
	
	CLB_6_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(139 downto 136),
	           snap_out     => CLB_6_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4619 downto 4488),
	           inputs       => CLB_6_5_inputs,
	           outputs      => CLB_6_5_outputs);
	
	CLB_6_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(143 downto 140),
	           snap_out     => CLB_6_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4751 downto 4620),
	           inputs       => CLB_6_6_inputs,
	           outputs      => CLB_6_6_outputs);
	
	CLB_7_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(147 downto 144),
	           snap_out     => CLB_7_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(4883 downto 4752),
	           inputs       => CLB_7_1_inputs,
	           outputs      => CLB_7_1_outputs);
	
	CLB_7_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(151 downto 148),
	           snap_out     => CLB_7_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5015 downto 4884),
	           inputs       => CLB_7_2_inputs,
	           outputs      => CLB_7_2_outputs);
	
	CLB_7_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(155 downto 152),
	           snap_out     => CLB_7_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5147 downto 5016),
	           inputs       => CLB_7_3_inputs,
	           outputs      => CLB_7_3_outputs);
	
	CLB_7_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(159 downto 156),
	           snap_out     => CLB_7_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5279 downto 5148),
	           inputs       => CLB_7_4_inputs,
	           outputs      => CLB_7_4_outputs);
	
	CLB_7_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(163 downto 160),
	           snap_out     => CLB_7_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5411 downto 5280),
	           inputs       => CLB_7_5_inputs,
	           outputs      => CLB_7_5_outputs);
	
	CLB_7_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(167 downto 164),
	           snap_out     => CLB_7_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5543 downto 5412),
	           inputs       => CLB_7_6_inputs,
	           outputs      => CLB_7_6_outputs);
	
	CLB_8_1: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(171 downto 168),
	           snap_out     => CLB_8_1_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5675 downto 5544),
	           inputs       => CLB_8_1_inputs,
	           outputs      => CLB_8_1_outputs);
	
	CLB_8_2: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(175 downto 172),
	           snap_out     => CLB_8_2_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5807 downto 5676),
	           inputs       => CLB_8_2_inputs,
	           outputs      => CLB_8_2_outputs);
	
	CLB_8_3: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(179 downto 176),
	           snap_out     => CLB_8_3_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(5939 downto 5808),
	           inputs       => CLB_8_3_inputs,
	           outputs      => CLB_8_3_outputs);
	
	CLB_8_4: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(183 downto 180),
	           snap_out     => CLB_8_4_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(6071 downto 5940),
	           inputs       => CLB_8_4_inputs,
	           outputs      => CLB_8_4_outputs);
	
	CLB_8_5: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(187 downto 184),
	           snap_out     => CLB_8_5_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(6203 downto 6072),
	           inputs       => CLB_8_5_inputs,
	           outputs      => CLB_8_5_outputs);
	
	CLB_8_6: entity work.CLB_clb_N4K4I10O4
	port map ( clk          => clk,
	           rst          => rst,
	           clk_app      => clk_app,
	           snap_in      => snap_in(191 downto 188),
	           snap_out     => CLB_8_6_snapshot_out,
	           snap_restore => snap_restore,
	           config       => config(6335 downto 6204),
	           inputs       => CLB_8_6_inputs,
	           outputs      => CLB_8_6_outputs);
	

end RTL;


--------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_wrapper is
	port ( clk          : in  std_ulogic;
	       rst          : in  std_ulogic;
	       --------------------------------------------------
	       clk_app      : in  std_ulogic;
	       rst_app      : in  std_ulogic;
	       snap_save    : in  std_ulogic;
	       snap_restore : in  std_ulogic;
	       --------------------------------------------------
               -- PGS 20190215 - Export shifted out config, so that we can
               -- freeze the VFPGA
	       config_out    : out  std_ulogic_vector(31 downto 0);
	       config_in    : in  std_ulogic_vector(31 downto 0);
	       config_valid : in  std_ulogic;
	       --------------------------------------------------
	       snap_in      : in  std_ulogic_vector(31 downto 0);
	       snap_out     : out std_ulogic_vector(31 downto 0);
	       snap_shift   : in  std_ulogic;
	       --------------------------------------------------
	       inputs       : in  std_ulogic_vector(55 downto 0);
	       outputs      : out std_ulogic_vector(55 downto 0));
end ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_wrapper;


architecture RTL of ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_wrapper is

	signal vFPGA_rst            : std_ulogic;
	signal vFPGA_config         : std_ulogic_vector(10951 downto 0) := (others => '0');
	signal vFPGA_snapshot_in    : std_ulogic_vector(191 downto 0) := (others => '0');
	signal vFPGA_snapshot_out   : std_ulogic_vector(191 downto 0) := (others => '0');
	signal vFPGA_inputs         : std_ulogic_vector(55 downto 0) := (others => '0');
	signal vFPGA_outputs        : std_ulogic_vector(55 downto 0) := (others => '0');
	signal vFPGA_outputs_registered : std_ulogic_vector(55 downto 0) := (others => '0');
                                
	signal config               : std_ulogic_vector(11623 downto 0) := (others => '0');
	signal snapshot             : std_ulogic_vector(191 downto 0) := (others => '0');
                                
	signal old_config_valid     : std_ulogic := '0';
	signal old_snap_shift       : std_ulogic := '0';
	signal old_snap_save        : std_ulogic := '0';

	signal io_reordering_config : std_ulogic_vector(671 downto 0) := (others => '0');
	signal input_choices        : std_ulogic_vector(63 downto 0) := (others => '0');
	signal output_choices       : std_ulogic_vector(63 downto 0) := (others => '0');

begin

	process (clk)
	begin
		if rising_edge(clk) then
			vFPGA_rst <= rst or rst_app;
		end if;
	end process;


	vFPGA_matrix: entity work.ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_matrix
	port map ( clk          => clk,
	           rst          => vFPGA_rst,
	           clk_app      => clk_app,
	           config       => vFPGA_config,
	           snap_in      => vFPGA_snapshot_in,
	           snap_out     => vFPGA_snapshot_out,
	           snap_restore => snap_restore,
	           inputs       => vFPGA_inputs,
	           outputs      => vFPGA_outputs);


	io_reordering_config <= config(11623 downto 10952);
	vFPGA_config <= config(10951 downto 0);


	process (clk)
	begin
		if rising_edge(clk) then
			old_config_valid <= config_valid;
			if config_valid = '1' and old_config_valid = '0' then
                                config(11623 downto 11592) <= config_in;
				config(11591 downto 0) <= config(11623 downto 32);
                                -- PGS 20190215: Allow reading back of config
                                -- as well, to make freezing possible.
                                -- We output the word that will be shifted out
                                -- next time, so that we can see the first word
                                -- of config after the last has been loaded, so
                                -- that it is possible to read and write the
                                -- config in a continuous loop.
                                config_out <= config(63 downto 32);
			end if;
		end if;
	end process;


	process (clk)
	begin
		if rising_edge(clk) then
			old_snap_shift <= snap_shift;
			old_snap_save <= snap_save;
			if snap_save = '1' and old_snap_save = '0' then
				snapshot(191 downto 0) <= vFPGA_snapshot_out;
			elsif snap_shift = '1' and old_snap_shift = '0' then
				snapshot(191 downto 160) <= snap_in;
				snapshot(159 downto 0) <= snapshot(191 downto 32);
			end if;
		end if;
	end process;
	snap_out <= snapshot(31 downto 0);

	vFPGA_snapshot_in <= snapshot(191 downto 0);


	input_choices <= "00000000" & inputs;
	output_choices <= "00000000" & vFPGA_outputs_registered;

	process (clk)
	begin
		if rising_edge(clk) then
			-- INPUTS --
			vFPGA_inputs(0) <= input_choices(to_integer(unsigned(io_reordering_config(5 downto 0))));
			vFPGA_inputs(1) <= input_choices(to_integer(unsigned(io_reordering_config(11 downto 6))));
			vFPGA_inputs(2) <= input_choices(to_integer(unsigned(io_reordering_config(17 downto 12))));
			vFPGA_inputs(3) <= input_choices(to_integer(unsigned(io_reordering_config(23 downto 18))));
			vFPGA_inputs(4) <= input_choices(to_integer(unsigned(io_reordering_config(29 downto 24))));
			vFPGA_inputs(5) <= input_choices(to_integer(unsigned(io_reordering_config(35 downto 30))));
			vFPGA_inputs(6) <= input_choices(to_integer(unsigned(io_reordering_config(41 downto 36))));
			vFPGA_inputs(7) <= input_choices(to_integer(unsigned(io_reordering_config(47 downto 42))));
			vFPGA_inputs(8) <= input_choices(to_integer(unsigned(io_reordering_config(53 downto 48))));
			vFPGA_inputs(9) <= input_choices(to_integer(unsigned(io_reordering_config(59 downto 54))));
			vFPGA_inputs(10) <= input_choices(to_integer(unsigned(io_reordering_config(65 downto 60))));
			vFPGA_inputs(11) <= input_choices(to_integer(unsigned(io_reordering_config(71 downto 66))));
			vFPGA_inputs(12) <= input_choices(to_integer(unsigned(io_reordering_config(77 downto 72))));
			vFPGA_inputs(13) <= input_choices(to_integer(unsigned(io_reordering_config(83 downto 78))));
			vFPGA_inputs(14) <= input_choices(to_integer(unsigned(io_reordering_config(89 downto 84))));
			vFPGA_inputs(15) <= input_choices(to_integer(unsigned(io_reordering_config(95 downto 90))));
			vFPGA_inputs(16) <= input_choices(to_integer(unsigned(io_reordering_config(101 downto 96))));
			vFPGA_inputs(17) <= input_choices(to_integer(unsigned(io_reordering_config(107 downto 102))));
			vFPGA_inputs(18) <= input_choices(to_integer(unsigned(io_reordering_config(113 downto 108))));
			vFPGA_inputs(19) <= input_choices(to_integer(unsigned(io_reordering_config(119 downto 114))));
			vFPGA_inputs(20) <= input_choices(to_integer(unsigned(io_reordering_config(125 downto 120))));
			vFPGA_inputs(21) <= input_choices(to_integer(unsigned(io_reordering_config(131 downto 126))));
			vFPGA_inputs(22) <= input_choices(to_integer(unsigned(io_reordering_config(137 downto 132))));
			vFPGA_inputs(23) <= input_choices(to_integer(unsigned(io_reordering_config(143 downto 138))));
			vFPGA_inputs(24) <= input_choices(to_integer(unsigned(io_reordering_config(149 downto 144))));
			vFPGA_inputs(25) <= input_choices(to_integer(unsigned(io_reordering_config(155 downto 150))));
			vFPGA_inputs(26) <= input_choices(to_integer(unsigned(io_reordering_config(161 downto 156))));
			vFPGA_inputs(27) <= input_choices(to_integer(unsigned(io_reordering_config(167 downto 162))));
			vFPGA_inputs(28) <= input_choices(to_integer(unsigned(io_reordering_config(173 downto 168))));
			vFPGA_inputs(29) <= input_choices(to_integer(unsigned(io_reordering_config(179 downto 174))));
			vFPGA_inputs(30) <= input_choices(to_integer(unsigned(io_reordering_config(185 downto 180))));
			vFPGA_inputs(31) <= input_choices(to_integer(unsigned(io_reordering_config(191 downto 186))));
			vFPGA_inputs(32) <= input_choices(to_integer(unsigned(io_reordering_config(197 downto 192))));
			vFPGA_inputs(33) <= input_choices(to_integer(unsigned(io_reordering_config(203 downto 198))));
			vFPGA_inputs(34) <= input_choices(to_integer(unsigned(io_reordering_config(209 downto 204))));
			vFPGA_inputs(35) <= input_choices(to_integer(unsigned(io_reordering_config(215 downto 210))));
			vFPGA_inputs(36) <= input_choices(to_integer(unsigned(io_reordering_config(221 downto 216))));
			vFPGA_inputs(37) <= input_choices(to_integer(unsigned(io_reordering_config(227 downto 222))));
			vFPGA_inputs(38) <= input_choices(to_integer(unsigned(io_reordering_config(233 downto 228))));
			vFPGA_inputs(39) <= input_choices(to_integer(unsigned(io_reordering_config(239 downto 234))));
			vFPGA_inputs(40) <= input_choices(to_integer(unsigned(io_reordering_config(245 downto 240))));
			vFPGA_inputs(41) <= input_choices(to_integer(unsigned(io_reordering_config(251 downto 246))));
			vFPGA_inputs(42) <= input_choices(to_integer(unsigned(io_reordering_config(257 downto 252))));
			vFPGA_inputs(43) <= input_choices(to_integer(unsigned(io_reordering_config(263 downto 258))));
			vFPGA_inputs(44) <= input_choices(to_integer(unsigned(io_reordering_config(269 downto 264))));
			vFPGA_inputs(45) <= input_choices(to_integer(unsigned(io_reordering_config(275 downto 270))));
			vFPGA_inputs(46) <= input_choices(to_integer(unsigned(io_reordering_config(281 downto 276))));
			vFPGA_inputs(47) <= input_choices(to_integer(unsigned(io_reordering_config(287 downto 282))));
			vFPGA_inputs(48) <= input_choices(to_integer(unsigned(io_reordering_config(293 downto 288))));
			vFPGA_inputs(49) <= input_choices(to_integer(unsigned(io_reordering_config(299 downto 294))));
			vFPGA_inputs(50) <= input_choices(to_integer(unsigned(io_reordering_config(305 downto 300))));
			vFPGA_inputs(51) <= input_choices(to_integer(unsigned(io_reordering_config(311 downto 306))));
			vFPGA_inputs(52) <= input_choices(to_integer(unsigned(io_reordering_config(317 downto 312))));
			vFPGA_inputs(53) <= input_choices(to_integer(unsigned(io_reordering_config(323 downto 318))));
			vFPGA_inputs(54) <= input_choices(to_integer(unsigned(io_reordering_config(329 downto 324))));
			vFPGA_inputs(55) <= input_choices(to_integer(unsigned(io_reordering_config(335 downto 330))));
			-- OUTPUTS --
			vFPGA_outputs_registered <= vFPGA_outputs;
			outputs(0) <= output_choices(to_integer(unsigned(io_reordering_config(341 downto 336))));
			outputs(1) <= output_choices(to_integer(unsigned(io_reordering_config(347 downto 342))));
			outputs(2) <= output_choices(to_integer(unsigned(io_reordering_config(353 downto 348))));
			outputs(3) <= output_choices(to_integer(unsigned(io_reordering_config(359 downto 354))));
			outputs(4) <= output_choices(to_integer(unsigned(io_reordering_config(365 downto 360))));
			outputs(5) <= output_choices(to_integer(unsigned(io_reordering_config(371 downto 366))));
			outputs(6) <= output_choices(to_integer(unsigned(io_reordering_config(377 downto 372))));
			outputs(7) <= output_choices(to_integer(unsigned(io_reordering_config(383 downto 378))));
			outputs(8) <= output_choices(to_integer(unsigned(io_reordering_config(389 downto 384))));
			outputs(9) <= output_choices(to_integer(unsigned(io_reordering_config(395 downto 390))));
			outputs(10) <= output_choices(to_integer(unsigned(io_reordering_config(401 downto 396))));
			outputs(11) <= output_choices(to_integer(unsigned(io_reordering_config(407 downto 402))));
			outputs(12) <= output_choices(to_integer(unsigned(io_reordering_config(413 downto 408))));
			outputs(13) <= output_choices(to_integer(unsigned(io_reordering_config(419 downto 414))));
			outputs(14) <= output_choices(to_integer(unsigned(io_reordering_config(425 downto 420))));
			outputs(15) <= output_choices(to_integer(unsigned(io_reordering_config(431 downto 426))));
			outputs(16) <= output_choices(to_integer(unsigned(io_reordering_config(437 downto 432))));
			outputs(17) <= output_choices(to_integer(unsigned(io_reordering_config(443 downto 438))));
			outputs(18) <= output_choices(to_integer(unsigned(io_reordering_config(449 downto 444))));
			outputs(19) <= output_choices(to_integer(unsigned(io_reordering_config(455 downto 450))));
			outputs(20) <= output_choices(to_integer(unsigned(io_reordering_config(461 downto 456))));
			outputs(21) <= output_choices(to_integer(unsigned(io_reordering_config(467 downto 462))));
			outputs(22) <= output_choices(to_integer(unsigned(io_reordering_config(473 downto 468))));
			outputs(23) <= output_choices(to_integer(unsigned(io_reordering_config(479 downto 474))));
			outputs(24) <= output_choices(to_integer(unsigned(io_reordering_config(485 downto 480))));
			outputs(25) <= output_choices(to_integer(unsigned(io_reordering_config(491 downto 486))));
			outputs(26) <= output_choices(to_integer(unsigned(io_reordering_config(497 downto 492))));
			outputs(27) <= output_choices(to_integer(unsigned(io_reordering_config(503 downto 498))));
			outputs(28) <= output_choices(to_integer(unsigned(io_reordering_config(509 downto 504))));
			outputs(29) <= output_choices(to_integer(unsigned(io_reordering_config(515 downto 510))));
			outputs(30) <= output_choices(to_integer(unsigned(io_reordering_config(521 downto 516))));
			outputs(31) <= output_choices(to_integer(unsigned(io_reordering_config(527 downto 522))));
			outputs(32) <= output_choices(to_integer(unsigned(io_reordering_config(533 downto 528))));
			outputs(33) <= output_choices(to_integer(unsigned(io_reordering_config(539 downto 534))));
			outputs(34) <= output_choices(to_integer(unsigned(io_reordering_config(545 downto 540))));
			outputs(35) <= output_choices(to_integer(unsigned(io_reordering_config(551 downto 546))));
			outputs(36) <= output_choices(to_integer(unsigned(io_reordering_config(557 downto 552))));
			outputs(37) <= output_choices(to_integer(unsigned(io_reordering_config(563 downto 558))));
			outputs(38) <= output_choices(to_integer(unsigned(io_reordering_config(569 downto 564))));
			outputs(39) <= output_choices(to_integer(unsigned(io_reordering_config(575 downto 570))));
			outputs(40) <= output_choices(to_integer(unsigned(io_reordering_config(581 downto 576))));
			outputs(41) <= output_choices(to_integer(unsigned(io_reordering_config(587 downto 582))));
			outputs(42) <= output_choices(to_integer(unsigned(io_reordering_config(593 downto 588))));
			outputs(43) <= output_choices(to_integer(unsigned(io_reordering_config(599 downto 594))));
			outputs(44) <= output_choices(to_integer(unsigned(io_reordering_config(605 downto 600))));
			outputs(45) <= output_choices(to_integer(unsigned(io_reordering_config(611 downto 606))));
			outputs(46) <= output_choices(to_integer(unsigned(io_reordering_config(617 downto 612))));
			outputs(47) <= output_choices(to_integer(unsigned(io_reordering_config(623 downto 618))));
			outputs(48) <= output_choices(to_integer(unsigned(io_reordering_config(629 downto 624))));
			outputs(49) <= output_choices(to_integer(unsigned(io_reordering_config(635 downto 630))));
			outputs(50) <= output_choices(to_integer(unsigned(io_reordering_config(641 downto 636))));
			outputs(51) <= output_choices(to_integer(unsigned(io_reordering_config(647 downto 642))));
			outputs(52) <= output_choices(to_integer(unsigned(io_reordering_config(653 downto 648))));
			outputs(53) <= output_choices(to_integer(unsigned(io_reordering_config(659 downto 654))));
			outputs(54) <= output_choices(to_integer(unsigned(io_reordering_config(665 downto 660))));
			outputs(55) <= output_choices(to_integer(unsigned(io_reordering_config(671 downto 666))));
		end if;
	end process;

end RTL;

--------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity vFPGA_clock_controler is
	port (clk               : in  std_ulogic;
	      rst               : in  std_ulogic;
	      clk_div           : in  std_ulogic_vector(9 downto 0);  -- How much to divide the physical clock to get the virtual clock (the actual value will be one more than the one written)
	      clk_cont_in       : in  std_ulogic_vector(23 downto 0); -- How many virtual clock cycles you want, 0 -> stoped, 111..1 -> never stop
	      clk_cont_in_valid : in  std_ulogic;
	      continue_clk_app  : in  std_ulogic;
	      clk_cont_out      : out std_ulogic_vector(23 downto 0); -- The remaining clock cycles
		  done              : out std_ulogic;                     -- Is set to one when the virtual clock is stoped (clk_count_out == 0)
		  clk_app           : out std_ulogic);                    -- The virtual clock, active for one physical clock cycle
end vFPGA_clock_controler;


architecture Behavioral of vFPGA_clock_controler is

	signal clk_div_counter   : std_ulogic_vector(9 downto 0) := (others => '0');
	signal clk_cycle_counter : std_ulogic_vector(23 downto 0) := (others => '0');
	signal clk_div_counter_down : std_ulogic_vector(9 downto 0) := (others => '0');

begin

	-- Virtual clock is active during only one physical clock cycle --
	process (clk)
	begin
		if rising_edge(clk) then
			if clk_div_counter = "0000000000" then
				clk_app <= '1';
			else
				clk_app <= '0';
			end if;
		end if;
	end process;


	-- Divisor counter --
	clk_div_counter_down <= std_ulogic_vector(unsigned(clk_div_counter) - 1);
	process (clk)
	begin
		if rising_edge(clk) then
			if continue_clk_app = '1' then
				if clk_div_counter = "0000000000" then
					clk_div_counter <= clk_div;
				else
					clk_div_counter <= clk_div_counter_down;
				end if;
			elsif clk_cycle_counter = x"000000" or rst = '1' or clk_div_counter = "0000000000" or clk_cont_in_valid = '1' then
				clk_div_counter <= clk_div;
			else
				clk_div_counter <= clk_div_counter_down;
			end if;
		end if;
	end process;


	-- Cycle counter --
	process (clk)
	begin
		if rising_edge(clk) then
			if rst = '1' then
				clk_cycle_counter <= x"000000";
			elsif clk_cont_in_valid = '1' then
				clk_cycle_counter <= clk_cont_in;
			elsif clk_div_counter = "0000000000" and clk_cycle_counter /= x"000000" and clk_cycle_counter /= x"ffffff" then
				clk_cycle_counter <= std_ulogic_vector(unsigned(clk_cycle_counter) - 1);
			end if;
		end if;
	end process;
				
	clk_cont_out <= clk_cycle_counter;


	-- done --
	process(clk)
	begin
		if rising_edge(clk) then
			if clk_cycle_counter = x"000000" then
				done <= '1';
			else
				done <= '0';
			end if;
		end if;
	end process;

end Behavioral;


--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- 00 pres 1
-- 04 pres 2
-- 08 pres 3
-- 0c SR
-- 10 CR
-- 14 DMAINADDRS
-- 18 DMAINADDRE
-- 1c DMAOUTADDRS
-- 20 DMAOUTADDRE
-- 24 MEMADDROFFSET
-- 28 CLKDIV
-- 2c CLKCNT
-- 30 CONFIG
-- 34 SNAPIN
-- 38 SNAPOUT

entity VFPGA_WRAPPER is
	Port ( -- WISHBONE --------------------------------------------
		   CLK_I          : in  std_logic;                     
		   RST_I          : in  std_logic;                     
		   -- WISHBONE SLAVE INTERFACE ----------------------------
		   SLAVE_CYC_I    : in  std_logic;                     
		   SLAVE_STB_I    : in  std_logic;                     
		   SLAVE_WE_I     : in  std_logic;                     
		   SLAVE_SEL_I    : in  std_logic_vector(3 downto 0);  
		   SLAVE_ADR_I    : in  std_logic_vector(7 downto 0); 
		   SLAVE_DAT_I    : in  std_logic_vector(31 downto 0); 
		   SLAVE_DAT_O    : out std_logic_vector(31 downto 0); 
		   SLAVE_ACK_O    : out std_logic;
		   --------------------------------------------------------
   	 	   VFPGA_CLK      : out std_logic;	
           INPUTS         : in  std_logic_vector(55 downto 0);
           OUTPUTS        : out std_logic_vector(55 downto 0));
end VFPGA_WRAPPER;


architecture Behavioral of VFPGA_WRAPPER is

	signal CLK_I_u          : std_ulogic := '0';
	signal RST_I_u          : std_ulogic := '0';
	signal SLAVE_CYC_I_u    : std_ulogic := '0';
	signal SLAVE_STB_I_u    : std_ulogic := '0';
	signal SLAVE_WE_I_u     : std_ulogic := '0';
	signal SLAVE_SEL_I_u    : std_ulogic_vector(3 downto 0) := (others => '0');  
	signal SLAVE_ADR_I_u    : std_ulogic_vector(7 downto 0) := (others => '0'); 
	signal SLAVE_DAT_I_u    : std_ulogic_vector(31 downto 0) := (others => '0'); 
	signal SLAVE_DAT_O_u    : std_ulogic_vector(31 downto 0) := (others => '0'); 
	signal SLAVE_ACK_O_u    : std_ulogic := '0';
	signal MASTER_CYC_O_u   : std_ulogic := '0';
    signal MASTER_STB_O_u   : std_ulogic := '0';
    signal MASTER_WE_O_u    : std_ulogic := '0';
    signal MASTER_SEL_O_u   : std_ulogic_vector(3 downto 0) := (others => '0');
    signal MASTER_ADR_O_u   : std_ulogic_vector(29 downto 0) := (others => '0');
    signal MASTER_DAT_O_u   : std_ulogic_vector(31 downto 0) := (others => '0');
    signal MASTER_DAT_I_u   : std_ulogic_vector(31 downto 0) := (others => '0');
    signal MASTER_ACK_I_u   : std_ulogic := '0';
	signal INTERRUPT_u      : std_ulogic := '0';
                                   
	signal clk_app                 : std_ulogic := '0';
	signal vFPGA_snap_save         : std_ulogic := '0';
	signal vFPGA_snap_restore      : std_ulogic := '0';
	signal vFPGA_snap_in           : std_ulogic_vector(31 downto 0) := (others => '0');
	signal vFPGA_snap_out          : std_ulogic_vector(31 downto 0) := (others => '0');
	signal vFPGA_snap_shift        : std_ulogic := '0';
	signal vFPGA_config_in         : std_ulogic_vector(31 downto 0) := (others => '0');
	signal vFPGA_config_valid      : std_ulogic := '0';
	signal vFPGA_inputs            : std_ulogic_vector(55 downto 0) := (others => '0');
	signal vFPGA_outputs           : std_ulogic_vector(55 downto 0) := (others => '0');
	signal clk_done_IE             : std_logic := '0';

	signal reg_rst_app             : std_ulogic := '0';
	signal reg_clk_div             : std_ulogic_vector(9 downto 0) := (others => '0');
	signal reg_clk_cycle_counter   : std_ulogic_vector(23 downto 0) := (others => '0');

	signal clk_cycle_counter_valid : std_ulogic := '0';

	signal clk_cycle_counter_remainder : std_ulogic_vector(23 downto 0) := (others => '0');
	signal clk_cycle_counter_done  : std_ulogic := '0';

	signal global_interrupt        : std_ulogic := '0';
	signal global_interrupt_IE     : std_ulogic := '0';

	signal write_config            : std_ulogic := '0';
	signal old_write_config        : std_ulogic := '0';

	signal write_snap_in           : std_ulogic := '0';
	signal read_snap_out           : std_ulogic := '0';
	signal old_write_snap_in       : std_ulogic := '0';
	signal old_read_snap_out       : std_ulogic := '0';

	signal write_snap_save         : std_ulogic := '0';
	signal write_snap_restore      : std_ulogic := '0';
	signal old_write_snap_save     : std_ulogic := '0';
	signal old_write_snap_restore  : std_ulogic := '0';

	signal write_clkcnt            : std_ulogic := '0';
	signal old_write_clkcnt        : std_ulogic := '0';

begin

	CLK_I_u        <= std_ulogic(CLK_I);
	RST_I_u        <= std_ulogic(RST_I);
	SLAVE_CYC_I_u  <= std_ulogic(SLAVE_CYC_I);
	SLAVE_STB_I_u  <= std_ulogic(SLAVE_STB_I);
	SLAVE_WE_I_u   <= std_ulogic(SLAVE_WE_I);
	SLAVE_SEL_I_u  <= std_ulogic_vector(SLAVE_SEL_I);
	SLAVE_ADR_I_u  <= std_ulogic_vector(SLAVE_ADR_I);
	SLAVE_DAT_I_u  <= std_ulogic_vector(SLAVE_DAT_I);

	SLAVE_DAT_O    <= std_logic_vector(SLAVE_DAT_O_u);
	SLAVE_ACK_O    <= std_logic(SLAVE_ACK_O_u);

	VFPGA_CLK      <= std_logic(clk_app);

	process (CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			if RST_I_u = '1' then
				INTERRUPT_u <= '0';
				global_interrupt <= '0';
			else
				INTERRUPT_u <= global_interrupt and global_interrupt_IE;
				global_interrupt <= (clk_cycle_counter_done and clk_done_IE);
			end if;
		end if;
	end process;


	vFPGA: entity work.ARCH8X6W16N4I10K4FCI4FCO8PFI8PFO8IOPB2_wrapper
	port map ( clk          => CLK_I_u,
	           rst          => RST_I_u,
	           clk_app      => clk_app,
	           rst_app      => reg_rst_app,
	           snap_save    => vFPGA_snap_save,
	           snap_restore => vFPGA_snap_restore,
	           config_in    => vFPGA_config_in,
	           config_valid => vFPGA_config_valid,
	           snap_in      => vFPGA_snap_in,
	           snap_out     => vFPGA_snap_out,
	           snap_shift   => vFPGA_snap_shift,
	           inputs       => vFPGA_inputs,
	           outputs      => vFPGA_outputs);


	CLK_CTRL: entity work.vFPGA_clock_controler
	port map ( clk               => CLK_I_u,
	           rst               => RST_I_u,
	           clk_div           => reg_clk_div,
	           clk_cont_in       => reg_clk_cycle_counter,
	           clk_cont_in_valid => clk_cycle_counter_valid,
	           continue_clk_app  => '0',
	           clk_cont_out      => clk_cycle_counter_remainder,
		       done              => clk_cycle_counter_done,
		       clk_app           => clk_app);


	-- Read process --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			SLAVE_DAT_O_u <= (others => '0');
			if (RST_I_u = '0') and (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') then
				SLAVE_DAT_O_u  <= (others => '0');
				case SLAVE_ADR_I_u is
					when "00000000" => -- PRES1
						SLAVE_DAT_O_u( 5 downto  0) <= "000111"; -- width
						SLAVE_DAT_O_u(11 downto  6) <= "000101"; -- height
						SLAVE_DAT_O_u(17 downto 12) <= "000111";  -- Logical wire cardinality (= W/2)
						SLAVE_DAT_O_u(21 downto 18) <= "0011";    -- N
						SLAVE_DAT_O_u(28 downto 22) <= "0001001";    -- I
						SLAVE_DAT_O_u(31 downto 29) <= "011";    -- K
					when "00000001" => -- PRES2
						SLAVE_DAT_O_u(22 downto  0) <= "00000000010110101101000"; -- Bitstream size in bits
						SLAVE_DAT_O_u(31 downto 23) <= "000111000"; -- Number of IO bits (= nb inputs = nb outputs)
					when "00000010" => -- PRES3
						SLAVE_DAT_O_u( 5 downto  0) <= "000000"; -- DMA word width
						SLAVE_DAT_O_u(11 downto  6) <= "000000"; -- MEM word width
						SLAVE_DAT_O_u(17 downto 12) <= "000000"; -- MEM address width
						SLAVE_DAT_O_u(18) <= '0'; -- With DMA ?
						SLAVE_DAT_O_u(19) <= '0'; -- With MEM access ?
						SLAVE_DAT_O_u(20) <= '0'; -- With interrupt pin ?
						SLAVE_DAT_O_u(31 downto 21) <= "10011001010"; -- Architecture file SHA1 11 LSB bits
					when "00000011" => -- SR
						SLAVE_DAT_O_u(5 downto  0) <= "110" & "0" & clk_cycle_counter_done & reg_rst_app;
						SLAVE_DAT_O_u(8) <= global_interrupt;
					when "00000100" => -- CR
						SLAVE_DAT_O_u(1 downto  0) <= '0' & reg_rst_app;
						SLAVE_DAT_O_u(8) <= global_interrupt_IE;
						SLAVE_DAT_O_u(12) <= clk_done_IE;
					when "00001010" => -- CLKDIV
						SLAVE_DAT_O_u(9 downto 0) <= reg_clk_div;
					when "00001011" => -- CLKCNT
						SLAVE_DAT_O_u(23 downto 0) <= clk_cycle_counter_remainder;
					when "00001100" => -- CONFIG
						SLAVE_DAT_O_u <= vFPGA_config_in;
					when "00001101" => -- SNAPIN
						SLAVE_DAT_O_u <= vFPGA_snap_in;
					when "00001110" => -- SNAPOUT
						SLAVE_DAT_O_u <= vFPGA_snap_out;
					when others =>
						null;
				end case;
			end if;
		end if;
	end process;


	-- Write control register --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			if RST_I_u = '1' then
				reg_rst_app <= '1';
				global_interrupt_IE <= '0';
				clk_done_IE <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00000100") then
				reg_rst_app <= SLAVE_DAT_I_u(0);
				global_interrupt_IE <= SLAVE_DAT_I_u(8);
				clk_done_IE <= SLAVE_DAT_I_u(12);
			end if;
		end if;
	end process;


	-- Snap save --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_write_snap_save  <= write_snap_save;
			vFPGA_snap_save <= write_snap_save and not (old_write_snap_save);
			if RST_I_u = '1' then
				write_snap_save <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00000100") and (SLAVE_SEL_I_u(0) = '1') and (SLAVE_DAT_I_u(2) = '1') then
				write_snap_save <= '1';
			else
				write_snap_save <= '0';
			end if;
		end if;
	end process;


	-- Snap restore --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_write_snap_restore <= write_snap_restore;
			vFPGA_snap_restore <= write_snap_restore and not (old_write_snap_restore);
			if RST_I_u = '1' then
				write_snap_restore <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00000100") and (SLAVE_SEL_I_u(0) = '1') and (SLAVE_DAT_I_u(3) = '1') then
				write_snap_restore <= '1';
			else
				write_snap_restore <= '0';
			end if;
		end if;
	end process;


	-- Write vclk divisor --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			if RST_I_u = '1' then
				reg_clk_div <= (others => '1');
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00001010") then
				reg_clk_div <= SLAVE_DAT_I_u(9 downto 0);
			end if;
		end if;
	end process;


	-- Write vclk cycle counter --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_write_clkcnt <= write_clkcnt;
			clk_cycle_counter_valid <= write_clkcnt and not(old_write_clkcnt);
			if RST_I_u = '1' then
				reg_clk_cycle_counter <= (others => '0');
				write_clkcnt <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00001011") then
				reg_clk_cycle_counter <= SLAVE_DAT_I_u(23 downto 0);
				write_clkcnt <= '1';
			else
				write_clkcnt <= '0';
			end if;
		end if;
	end process;


	-- Write vFPGA config word --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_write_config <= write_config;
			vFPGA_config_valid <= write_config and not(old_write_config);
			if RST_I_u = '1' then
				vFPGA_config_in <= (others => '0');
				write_config <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00001100") then
				vFPGA_config_in <= SLAVE_DAT_I_u;
				write_config <= '1';
			else
				write_config <= '0';
			end if;
		end if;
	end process;


	-- Write vFPGA snapshot word --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_write_snap_in <= write_snap_in;
			if RST_I_u = '1' then
				vFPGA_snap_in <= (others => '0');
				write_snap_in <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '1') and (SLAVE_ADR_I_u = "00001101") then
				vFPGA_snap_in <= SLAVE_DAT_I_u;
				write_snap_in <= '1';
			else
				write_snap_in <= '0';
			end if;
		end if;
	end process;


	-- Read vFPGA snapshot word --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			old_read_snap_out <= read_snap_out;
			if RST_I_u = '1' then
				read_snap_out <= '0';
			elsif (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_WE_I_u = '0') and (SLAVE_ADR_I_u = "00001110") then
				read_snap_out <= '1';
			else
				read_snap_out <= '0';
			end if;
		end if;
	end process;


	-- Shift snapshot when writting snapin and after reading snapout --
	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			vFPGA_snap_shift <= (write_snap_in and not(old_write_snap_in)) or (not(read_snap_out) and old_read_snap_out);
		end if;
	end process;


	vFPGA_inputs <= std_ulogic_vector(INPUTS);
	OUTPUTS <= std_logic_vector(vFPGA_outputs);














	process(CLK_I_u)
	begin
		if rising_edge(CLK_I_u) then
			if (RST_I_u = '0') and (SLAVE_CYC_I_u = '1') and (SLAVE_STB_I_u = '1') and (SLAVE_ACK_O_u = '0') then
				SLAVE_ACK_O_u <= '1';
			else 
				SLAVE_ACK_O_u <= '0';
			end if;
		end if;
	end process;

end Behavioral;
               


-- Full signature --
--
-- 4a4203081c002d6899400000

