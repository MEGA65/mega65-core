library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use STD.textio.all;
use work.debugtools.all;
use work.cputypes.all;

entity test_readcomp is
end entity;

architecture foo of test_readcomp is

  type CharFile is file of character;

  signal clock40mhz : std_logic := '1';
  signal clock80mhz : std_logic := '1';
  -- $51 = DD, $28 = HD, $14 = ED
  signal cycles_per_interval : unsigned(7 downto 0) := x"16";
  
  signal cycle_count : integer := 0;

  signal gap_valid_in : std_logic := '0';
  signal gap_length_in : unsigned(15 downto 0) := (others => '0');
    
  signal gap_valid_out : std_logic := '0';
  signal gap_length_out : unsigned(15 downto 0) := (others => '0');

  signal gap_num : integer := 0;
  type gaps_t is array(0 to 10000) of integer;
  signal gap_lengths : gaps_t := (
22, 22, 22, 22, 22, 22, 23, 27, 35, 35, 44, 35, 35, 24, 57, 24, 
23, 56, 21, 24, 57, 22, 24, 28, 29, 36, 35, 25, 29, 23, 21, 22, 
22, 22, 22, 21, 22, 22, 23, 34, 21, 21, 23, 34, 24, 35, 29, 28, 
22, 23, 36, 35, 25, 44, 37, 36, 44, 36, 38, 44, 37, 36, 45, 36, 
37, 43, 36, 38, 45, 36, 37, 44, 36, 37, 45, 35, 37, 44, 36, 37, 
45, 34, 36, 44, 37, 37, 44, 36, 38, 44, 37, 36, 45, 36, 37, 43, 
36, 36, 46, 37, 37, 43, 36, 36, 45, 36, 37, 44, 37, 35, 44, 36, 
38, 45, 37, 36, 45, 36, 37, 44, 37, 33, 21, 21, 21, 22, 22, 22, 
22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 
22, 22, 22, 23, 21, 21, 21, 21, 21, 21, 23, 21, 21, 21, 21, 21, 
21, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 23, 22, 
22, 21, 22, 22, 22, 22, 22, 21, 21, 21, 23, 56, 21, 24, 57, 23, 
23, 55, 21, 23, 28, 34, 23, 57, 29, 36, 53, 30, 30, 49, 22, 22, 
22, 23, 26, 20, 22, 43, 27, 21, 23, 29, 42, 22, 22, 23, 50, 34, 
23, 34, 23, 33, 23, 28, 29, 51, 43, 24, 50, 35, 30, 42, 22, 23, 
28, 42, 42, 28, 43, 30, 44, 42, 23, 50, 35, 28, 23, 28, 36, 52, 
29, 36, 37, 44, 36, 30, 51, 29, 23, 24, 43, 29, 35, 24, 29, 30, 
43, 42, 28, 36, 52, 29, 30, 35, 24, 28, 29, 29, 31, 29, 24, 42, 
23, 26, 22, 34, 27, 23, 27, 23, 42, 23, 40, 28, 26, 22, 50, 41, 
22, 43, 50, 23, 36, 34, 22, 24, 35, 28, 27, 24, 29, 42, 22, 23, 
29, 34, 24, 27, 21, 22, 22, 24, 27, 23, 42, 22, 26, 22, 29, 35, 
28, 23, 23, 43, 41, 22, 50, 41, 22, 27, 23, 57, 58, 59, 35, 25, 
50, 23, 21, 22, 51, 42, 24, 50, 28, 36, 50, 24, 44, 42, 27, 22, 
24, 43, 50, 23, 43, 35, 36, 44, 30, 43, 36, 24, 24, 35, 35, 35, 
22, 23, 36, 44, 37, 36, 38, 45, 37, 29, 52, 35, 28, 28, 23, 33, 
23, 57, 35, 24, 35, 24, 28, 28, 23, 35, 30, 40, 27, 22, 29, 51, 
36, 30, 44, 43, 29, 37, 51, 31, 37, 28, 24, 27, 28, 58, 30, 29, 
29, 29, 24, 23, 23, 41, 21, 22, 50, 27, 22, 34, 24, 28, 22, 23, 
35, 34, 21, 22, 28, 42, 23, 23, 26, 22, 28, 23, 35, 49, 22, 21, 
22, 28, 29, 24, 29, 35, 25, 35, 25, 35, 27, 24, 29, 30, 29, 35, 
22, 23, 36, 51, 43, 25, 52, 44, 28, 22, 24, 34, 28, 50, 30, 35, 
42, 23, 23, 28, 43, 50, 42, 23, 42, 28, 43, 36, 37, 44, 29, 44, 
44, 29, 24, 41, 21, 23, 50, 41, 22, 28, 58, 28, 24, 29, 37, 59, 
59, 51, 30, 35, 43, 36, 37, 36, 44, 37, 35, 25, 59, 30, 51, 36, 
29, 30, 49, 22, 23, 42, 27, 22, 22, 24, 51, 34, 23, 28, 29, 51, 
36, 31, 46, 43, 30, 41, 22, 50, 35, 50, 29, 37, 30, 51, 30, 35, 
24, 28, 29, 37, 51, 29, 30, 28, 29, 29, 24, 36, 29, 24, 43, 24, 
28, 23, 43, 49, 23, 34, 28, 28, 24, 28, 34, 23, 27, 23, 41, 21, 
26, 21, 23, 42, 41, 22, 27, 22, 58, 35, 25, 51, 43, 24, 50, 23, 
43, 42, 48, 23, 42, 28, 43, 35, 34, 22, 23, 35, 37, 44, 36, 30, 
28, 24, 35, 24, 33, 22, 28, 42, 22, 23, 29, 43, 44, 29, 37, 28, 
23, 28, 28, 30, 28, 23, 22, 21, 22, 27, 23, 49, 33, 21, 23, 26, 
22, 27, 23, 34, 28, 28, 23, 28, 37, 28, 23, 27, 23, 33, 49, 42, 
27, 22, 23, 27, 36, 43, 51, 43, 23, 35, 37, 44, 28, 24, 42, 22, 
23, 28, 58, 58, 59, 43, 36, 37, 35, 25, 58, 30, 30, 49, 22, 22, 
24, 50, 50, 36, 31, 42, 23, 50, 35, 29, 51, 31, 37, 51, 29, 24, 
36, 29, 24, 44, 50, 23, 27, 35, 23, 27, 22, 23, 43, 57, 34, 23, 
49, 24, 44, 43, 29, 43, 36, 37, 44, 35, 24, 33, 23, 28, 44, 43, 
29, 29, 29, 28, 25, 52, 35, 23, 22, 23, 28, 27, 23, 26, 21, 35, 
51, 30, 36, 44, 37, 36, 43, 24, 29, 58, 45, 36, 37, 29, 30, 51, 
51, 36, 30, 36, 31, 52, 28, 24, 36, 28, 23, 28, 35, 24, 57, 35, 
25, 43, 29, 44, 35, 24, 35, 24, 28, 30, 29, 28, 24, 35, 30, 27, 
22, 22, 28, 36, 44, 25, 30, 57, 29, 30, 51, 36, 30, 50, 24, 29, 
36, 25, 43, 29, 44, 29, 29, 30, 28, 23, 23, 29, 36, 36, 30, 30, 
50, 23, 27, 34, 23, 28, 29, 29, 58, 30, 30, 43, 28, 29, 30, 44, 
30, 29, 29, 29, 23, 21, 20, 23, 22, 22, 22, 22, 23, 26, 21, 22, 
34, 21, 22, 22, 22, 22, 23, 27, 23, 33, 22, 22, 22, 22, 23, 28, 
27, 21, 23, 33, 26, 20, 22, 22, 24, 34, 22, 23, 27, 21, 21, 22, 
23, 28, 41, 22, 23, 28, 27, 22, 23, 41, 22, 26, 22, 34, 27, 23, 
21, 21, 22, 48, 21, 21, 22, 34, 23, 23, 35, 29, 28, 23, 27, 21, 
21, 22, 23, 28, 35, 24, 34, 24, 41, 20, 22, 28, 36, 29, 24, 29, 
29, 23, 24, 42, 28, 30, 35, 23, 23, 25, 27, 39, 27, 33, 49, 26, 
21, 21, 21, 22, 42, 22, 51, 49, 23, 22, 24, 42, 27, 21, 22, 34, 
22, 23, 35, 35, 30, 50, 29, 28, 24, 35, 30, 36, 43, 23, 22, 22, 
23, 27, 21, 22, 28, 43, 35, 24, 34, 25, 50, 41, 23, 41, 20, 22, 
29, 43, 30, 43, 36, 29, 24, 29, 37, 36, 44, 29, 24, 24, 43, 28, 
43, 43, 28, 29, 36, 25, 29, 24, 43, 22, 23, 27, 23, 40, 29, 50, 
42, 23, 34, 33, 21, 22, 29, 57, 29, 24, 22, 22, 23, 27, 23, 28, 
36, 42, 23, 50, 59, 58, 50, 23, 21, 22, 50, 29, 36, 44, 29, 23, 
24, 43, 36, 36, 36, 23, 24, 36, 38, 44, 37, 35, 29, 51, 35, 24, 
58, 30, 28, 25, 37, 30, 52, 34, 28, 35, 51, 30, 29, 50, 23, 22, 
22, 23, 27, 21, 23, 42, 26, 21, 22, 28, 42, 22, 22, 23, 51, 34, 
23, 33, 22, 33, 22, 28, 30, 51, 43, 24, 51, 36, 30, 42, 22, 23, 
28, 44, 44, 29, 45, 29, 44, 42, 23, 49, 34, 27, 23, 28, 36, 51, 
30, 36, 37, 44, 36, 30, 51, 29, 24, 24, 42, 27, 34, 22, 28, 29, 
46, 44, 30, 36, 51, 29, 30, 35, 24, 29, 29, 31, 30, 27, 23, 41, 
22, 27, 22, 34, 27, 23, 27, 23, 41, 23, 40, 28, 26, 22, 50, 41, 
22, 43, 50, 24, 35, 34, 21, 23, 34, 28, 29, 24, 29, 43, 22, 23, 
28, 34, 23, 27, 22, 22, 22, 24, 28, 23, 41, 21, 26, 21, 27, 35, 
28, 23, 23, 42, 41, 22, 50, 41, 23, 27, 23, 56, 58, 58, 35, 25, 
50, 23, 21, 23, 50, 41, 22, 49, 28, 35, 51, 25, 45, 42, 27, 21, 
23, 42, 48, 23, 43, 35, 36, 43, 30, 42, 33, 22, 23, 35, 36, 35, 
23, 24, 36, 43, 36, 37, 38, 44, 37, 29, 51, 36, 30, 28, 24, 34, 
23, 58, 36, 25, 35, 24, 29, 29, 24, 35, 29, 43, 23, 23, 28, 50, 
36, 30, 44, 43, 28, 37, 51, 30, 36, 28, 24, 28, 29, 58, 30, 29, 
30, 28, 23, 22, 23, 41, 21, 22, 50, 27, 24, 34, 23, 26, 20, 23, 
35, 34, 22, 23, 28, 42, 22, 23, 27, 22, 27, 23, 35, 49, 22, 21, 
23, 28, 28, 24, 28, 33, 22, 34, 23, 34, 29, 24, 29, 29, 30, 35, 
23, 22, 36, 51, 44, 25, 52, 43, 27, 21, 23, 34, 29, 50, 29, 37, 
43, 22, 23, 29, 44, 51, 42, 23, 43, 29, 44, 36, 37, 44, 30, 43, 
43, 27, 23, 41, 22, 23, 50, 42, 22, 28, 58, 28, 23, 28, 37, 58, 
60, 51, 30, 36, 44, 36, 37, 36, 46, 36, 37, 25, 59, 29, 52, 34, 
29, 29, 50, 22, 24, 43, 28, 22, 22, 24, 50, 35, 24, 29, 30, 50, 
36, 31, 44, 44, 30, 41, 22, 50, 36, 50, 29, 36, 32, 53, 31, 35, 
24, 29, 30, 36, 51, 29, 30, 28, 29, 29, 24, 36, 29, 25, 43, 24, 
27, 24, 44, 49, 23, 35, 29, 28, 23, 27, 33, 23, 27, 23, 41, 22, 
27, 20, 23, 42, 41, 23, 27, 22, 58, 35, 24, 51, 43, 23, 48, 23, 
42, 42, 48, 22, 41, 27, 43, 36, 36, 23, 23, 35, 37, 43, 36, 29, 
29, 25, 36, 25, 34, 22, 29, 43, 22, 24, 29, 44, 44, 30, 36, 29, 
24, 29, 29, 29, 29, 24, 23, 22, 23, 26, 22, 50, 34, 22, 23, 27, 
22, 27, 23, 34, 29, 28, 24, 29, 36, 29, 24, 28, 24, 36, 53, 43, 
28, 22, 22, 28, 36, 45, 51, 44, 25, 36, 37, 44, 28, 24, 42, 22, 
22, 28, 59, 58, 59, 43, 36, 37, 35, 25, 58, 29, 30, 49, 23, 22, 
23, 50, 51, 36, 31, 42, 23, 49, 34, 28, 51, 30, 37, 51, 28, 24, 
36, 28, 24, 44, 50, 24, 28, 34, 23, 27, 21, 22, 44, 57, 35,


                                  others => 0);
  
  
begin

  comp0: entity work.floppy_read_compensate port map (
    clock40mhz => clock40mhz,
    correction_enable => '1',
    cycles_per_interval => cycles_per_interval,
    gap_valid_in => gap_valid_in,
    gap_length_in => gap_length_in,
    gap_valid_out => gap_valid_out,
    gap_length_out => gap_length_out
    );
  
  process is
  begin
    while true loop
      clock40mhz <= '0';
      clock80mhz <= '0';
      wait for 5 ns;
      clock80mhz <= '1';
      wait for 5 ns;
      clock40mhz <= '1';
      clock80mhz <= '0';
      wait for 5 ns;
      clock80mhz <= '1';
      wait for 5 ns;
    end loop;
  end process;

  
  process (clock40mhz) is
  begin
    if rising_edge(clock40mhz) then      
 
      if cycle_count = 0 then
        cycle_count <= gap_lengths(gap_num)*3 - 1;
        gap_valid_in <= '1';
        gap_length_in <= to_unsigned(gap_lengths(gap_num)*3,16);
        gap_num <= gap_num + 1;
        if gap_lengths(gap_num) = 0 then
          assert false;
          gap_num <= 99999;
        end if;
      else
        cycle_count <= cycle_count - 1;
        gap_valid_in <= '0';
      end if;
      
    end if;
  end process;
  
end foo;
