module uart_rx_buffered (input clk, input [23:0] bit_rate_divisor, input UART_RX, output [7:0] data, output data_ready, input data_acknowledge);

endmodule
