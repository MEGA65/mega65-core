library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.debugtools.all;

--
entity charrom is
port (Clk : in std_logic;
        address : in integer range 0 to 4095;
        -- chip select, active low       
        cs : in std_logic;
        data_o : out std_logic_vector(7 downto 0);

        writeclk : in std_logic;
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        writecs : in std_logic;
        we : in std_logic;
        writeaddress : in unsigned(11 downto 0);
        data_i : in std_logic_vector(7 downto 0)
      );
end charrom;

architecture Behavioral of charrom is

-- 4K x 8bit pre-initialised RAM
-- Characters are from:
-- http://users.ices.utexas.edu/~lenharth/cs378/fall13/font8x8.h
-- Original copyright notice:
--  * 8x8 monochrome bitmap fonts for rendering
 --* Author: Daniel Hepper <daniel@hepper.net>
 --* 
 --* License: Public Domain
 --* 
 --* Based on:
 --* // Summary: font8x8.h
 --* // 8x8 monochrome bitmap fonts for rendering
 --* //
 --* // Author:
 --* //     Marcel Sondaar
 --* //     International Business Machines (public domain VGA fonts)
 --* //
 --* // License:
 --* //     Public Domain
 --* 
 --* Fetched from: http://dimensionalrift.homelinux.net/combuster/mos3/?p=viewsource&file=/modules/gfx/font8_8.asm

type ram_t is array (0 to 4095) of std_logic_vector(7 downto 0);
signal ram : ram_t := (
  x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

  -- and repeat 7 more times
  x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

    x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

    x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

    x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

    x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

    x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",

  x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",
  x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",
  x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",
  x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",
  x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",
  x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",
  x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",
  x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",
  x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",
  x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",
  x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",
  x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
  x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",
  x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",
  x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",
  x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",
  x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",
  x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",
  x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",
  x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",
  x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",
  x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",
  x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",
  x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",
  x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",
  x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",
  x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
  x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",
  x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",
  x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",
  x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",
  x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",
  x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",
  x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",
  x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",
  x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",
  x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",
  x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",
  x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",
  x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",
  x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",
  x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",
  x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",
  x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",
  x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",
  x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",
  x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",
  x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",
  x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",
  x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",
  x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00"
  
);

begin

--process for read and write operation.
PROCESS(Clk)
BEGIN
  --report "viciv reading charrom address $"
  --  & to_hstring(address)
  --  & " = " & integer'image(to_integer(address))
  --  & " -> $" & to_hstring(ram(to_integer(address)))
  --  severity note;
  data_o <= ram(address);          

  if(rising_edge(writeClk)) then 
    if writecs='1' then
      if(we='1') then
            ram(to_integer(writeaddress)) <= data_i;
      end if;
    end if;
  end if;
END PROCESS;

end Behavioral;
