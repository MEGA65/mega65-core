module uart_rx (input clk, input [15:0] bit_rate_divisor, input UART_RX, output [7:0] data, output data_ready, input data_acknowledge);

endmodule
