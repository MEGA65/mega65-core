library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-------------------------------------------------------------------------------

entity sid_tables is
	port (
          clock : in std_logic;
          sawtooth : in unsigned(11 downto 0);
          triangle : in unsigned(11 downto 0);
          st_out : out unsigned(7 downto 0) := x"00";
          p_t_out : out unsigned(7 downto 0) := x"00";
          ps_out : out unsigned(7 downto 0) := x"00";
          pst_out : out unsigned(7 downto 0) := x"00"
          );
end sid_tables;

architecture sequential of sid_tables is

  type array4k is array(0 to 4095) of unsigned(7 downto 0);

   signal table_st : array4k := (
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0e", x"0e", x"0e", x"0e", x"0f", x"0f", x"0f", x"0f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1e", x"1e", x"1f", x"1f", x"1f", x"1f", x"1f", x"1f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0e", x"0e", x"0e", x"0e", x"0f", x"0f", x"0f", x"1f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38"
     , x"3c", x"3c", x"3c", x"3c", x"3c", x"3c", x"3c", x"3e", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0e", x"0e", x"0e", x"0e", x"0f", x"0f", x"0f", x"0f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1c", x"1e", x"1e", x"1f", x"1f", x"1f", x"1f", x"3f", x"3f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0e", x"0e", x"0e", x"0e", x"0f", x"0f", x"1f", x"1f"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
     , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"83", x"83"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
     , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"87", x"87", x"87", x"8f"
     , x"c0", x"e0", x"e0", x"c0", x"c0", x"e0", x"e0", x"e0", x"e0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
     , x"c0", x"e0", x"e0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
     , x"c0", x"e0", x"e0", x"c0", x"c0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"c0", x"e0", x"c0", x"e0", x"e0"
     , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
     , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
     , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
     , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
     , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e3", x"e3"
     , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0"
     , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0"
     , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0"
     , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1"
     , x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8"
     , x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8"
     , x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc"
     , x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
  
  signal table_p_t : array4k := (
    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1c", x"00", x"3c", x"3f", x"3f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0c", x"5e", x"5f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"40", x"40", x"60", x"60", x"6f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"40"
    , x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"60", x"40", x"40", x"60", x"60", x"60", x"60", x"70", x"77"
    , x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"60", x"60", x"60"
    , x"40", x"40", x"40", x"60", x"60", x"60", x"60", x"70", x"60", x"60", x"60", x"70", x"70", x"70", x"78", x"7b"
    , x"60", x"60", x"60", x"70", x"60", x"70", x"70", x"70", x"70", x"70", x"70", x"78", x"78", x"78", x"78", x"7c"
    , x"78", x"78", x"78", x"7c", x"78", x"7c", x"7c", x"7e", x"7c", x"7e", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"8e", x"9f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"80", x"80", x"80"
    , x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"00", x"00", x"00", x"80", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"af"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a0", x"a0", x"a0", x"a0", x"b7"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"a0", x"a0", x"a0", x"a0", x"a0", x"b0", x"a0", x"b0", x"b0", x"bb"
    , x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"b0", x"b0", x"a0", x"b0", x"b0", x"b8", x"b0", x"b8", x"b8", x"bc"
    , x"b0", x"b8", x"b8", x"b8", x"b8", x"bc", x"bc", x"be", x"bc", x"bc", x"be", x"bf", x"be", x"bf", x"bf", x"bf"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"c0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"80", x"80", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"80", x"80", x"80", x"c0", x"80", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"cf"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"c0", x"c0", x"80", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d7"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d0", x"d0", x"d9"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d0", x"c0", x"d0", x"d0", x"d0", x"d0", x"d8", x"d8", x"dc"
    , x"d0", x"d0", x"d8", x"d8", x"d8", x"dc", x"dc", x"de", x"dc", x"dc", x"de", x"df", x"de", x"df", x"df", x"df"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"e0", x"e0", x"e0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"c0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e7"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e8"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e8", x"ec"
    , x"e0", x"e0", x"e0", x"e8", x"e8", x"e8", x"ec", x"ee", x"ec", x"ec", x"ec", x"ee", x"ee", x"ef", x"ef", x"ef"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"f0", x"f0", x"f0"
    , x"e0", x"e0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0"
    , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4"
    , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"f0", x"f4", x"f4", x"f6", x"f6", x"f7", x"f7", x"f7"
    , x"f0", x"f0", x"f0", x"f8", x"f0", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8"
    , x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fa", x"fa", x"fb", x"fb", x"fb"
    , x"f8", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fd", x"fd", x"fd"
    , x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
  
  signal table_ps : array4k := (
    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"1f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"0f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"17"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3b"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3d"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3e"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3f", x"00", x"0c", x"1c", x"3f", x"1e", x"3f", x"3f", x"3f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0b"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0a"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5e"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5f", x"00", x"00", x"00", x"5f", x"0c", x"5f", x"5f", x"5f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"47"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"43"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"65"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6e"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6f", x"00", x"40", x"40", x"6f", x"40", x"6f", x"6f", x"6f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"63"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"61"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"40", x"00", x"40", x"40", x"70"
    , x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"70", x"40", x"60", x"60", x"77", x"60", x"77", x"77", x"77"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"60", x"00", x"40", x"40", x"60", x"40", x"60", x"60", x"79"
    , x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"60", x"78"
    , x"40", x"60", x"60", x"60", x"60", x"60", x"60", x"78", x"60", x"70", x"70", x"78", x"70", x"79", x"7b", x"7b"
    , x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"70", x"60", x"60", x"60", x"70", x"60", x"70", x"70", x"7c"
    , x"60", x"70", x"70", x"70", x"70", x"70", x"70", x"7c", x"70", x"78", x"78", x"7c", x"78", x"7c", x"7c", x"7d"
    , x"70", x"78", x"78", x"78", x"78", x"78", x"78", x"7c", x"78", x"7c", x"7c", x"7e", x"7c", x"7e", x"7e", x"7e"
    , x"7c", x"7c", x"7c", x"7e", x"7e", x"7f", x"7f", x"7f", x"7e", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"ff"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"87"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"83"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"8d"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"00", x"80", x"80", x"8e"
    , x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"8f", x"80", x"80", x"80", x"9f", x"80", x"9f", x"9f", x"9f"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"00", x"80", x"80", x"87"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"83"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"81"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"84"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"87", x"80", x"80", x"80", x"87", x"80", x"8f", x"af", x"af"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80"
    , x"00", x"00", x"00", x"80", x"00", x"00", x"80", x"80", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"83"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"81"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a0", x"80", x"80", x"80", x"a0", x"80", x"a3", x"b7", x"b7"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"b1"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"b0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"b0", x"80", x"a0", x"a0", x"b0", x"a0", x"b8", x"b9", x"bb"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"a0", x"80", x"80", x"80", x"a0", x"80", x"a0", x"a0", x"b8"
    , x"80", x"a0", x"a0", x"a0", x"a0", x"a0", x"a0", x"b8", x"a0", x"b0", x"b0", x"b8", x"b0", x"bc", x"bc", x"bd"
    , x"a0", x"b0", x"b0", x"b0", x"b0", x"b8", x"b8", x"bc", x"b0", x"b8", x"b8", x"bc", x"b8", x"bc", x"be", x"be"
    , x"b8", x"bc", x"bc", x"be", x"bc", x"be", x"be", x"bf", x"be", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf"
    , x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80"
    , x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"81"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c7"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"c3"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"80", x"80", x"80", x"c0", x"80", x"c0", x"c0", x"c1"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"80", x"80", x"80", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c7", x"c0", x"c0", x"c0", x"c7", x"c0", x"cf", x"cf", x"cf"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"c0", x"80", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c3"
    , x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"c0", x"80", x"80", x"80", x"c0", x"80", x"c0", x"c0", x"c0"
    , x"80", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c1"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c1", x"c7", x"d7"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d0", x"c0", x"c0", x"c0", x"d0", x"c0", x"d0", x"d8", x"db"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d8"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"d8", x"c0", x"c0", x"c0", x"d8", x"d0", x"d8", x"d8", x"dd"
    , x"c0", x"c0", x"c0", x"d0", x"c0", x"d0", x"d0", x"dc", x"d0", x"d8", x"d8", x"dc", x"d8", x"dc", x"dc", x"de"
    , x"d8", x"dc", x"dc", x"de", x"dc", x"de", x"de", x"df", x"de", x"df", x"df", x"df", x"df", x"df", x"df", x"df"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e3"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"c0", x"c0", x"e0", x"c0", x"e0", x"e0", x"e1"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"c0", x"c0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"c0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e1", x"e3", x"e7"
    , x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"c0", x"e0", x"c0", x"c0", x"c0", x"e0", x"c0", x"e0", x"e0", x"e0"
    , x"c0", x"c0", x"c0", x"e0", x"c0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"eb"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e8", x"e0", x"e8", x"e8", x"ed"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"ec", x"e0", x"e0", x"e0", x"ec", x"e8", x"ec", x"ec", x"ee"
    , x"e8", x"e8", x"e8", x"ec", x"ec", x"ee", x"ee", x"ef", x"ec", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef", x"ef"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"f0"
    , x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"e0", x"f0", x"e0", x"e0", x"e0", x"f0", x"e0", x"f0", x"f0", x"f0"
    , x"e0", x"e0", x"e0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f3"
    , x"e0", x"e0", x"e0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0"
    , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f5"
    , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"f4", x"f6"
    , x"f0", x"f0", x"f0", x"f4", x"f0", x"f4", x"f6", x"f7", x"f4", x"f6", x"f6", x"f7", x"f7", x"f7", x"f7", x"f7"
    , x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f8", x"f8", x"f8"
    , x"f0", x"f0", x"f0", x"f8", x"f0", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f9"
    , x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fa"
    , x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fb", x"f8", x"fa", x"fa", x"fb", x"fb", x"fb", x"fb", x"fb"
    , x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc"
    , x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fd", x"fc", x"fc", x"fc", x"fd", x"fd", x"fd", x"fd", x"fd"
    , x"fc", x"fc", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe", x"fe"
    , x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
  
  
begin
  
  process (clock,sawtooth,triangle) is
  begin
    if rising_edge(clock) then
      st_out <= table_st(to_integer(sawtooth));
      p_t_out <= table_p_t(to_integer(triangle));
      ps_out <= table_ps(to_integer(sawtooth));
      
      if sawtooth < x"3ff" then   pst_out <= x"00";
      elsif sawtooth < x"400" then   pst_out <= x"1f";
      elsif sawtooth < x"7ee" then   pst_out <= x"00";
      elsif sawtooth < x"7ef" then   pst_out <= x"20";
      elsif sawtooth < x"7f0" then   pst_out <= x"70";
      elsif sawtooth < x"7f1" then   pst_out <= x"60";
      elsif sawtooth < x"7f2" then   pst_out <= x"20";
      elsif sawtooth < x"7f7" then   pst_out <= x"70";
      elsif sawtooth < x"7fa" then   pst_out <= x"78";
      elsif sawtooth < x"7fc" then   pst_out <= x"7c";
      elsif sawtooth < x"7fe" then   pst_out <= x"7e";
      elsif sawtooth < x"800" then   pst_out <= x"7f";
      elsif sawtooth < x"bfd" then   pst_out <= x"00";
      elsif sawtooth < x"bfe" then   pst_out <= x"08";
      elsif sawtooth < x"bff" then   pst_out <= x"1e";
      elsif sawtooth < x"c00" then   pst_out <= x"3f";
      elsif sawtooth < x"df7" then   pst_out <= x"00";
      elsif sawtooth < x"dfe" then   pst_out <= x"80";
      elsif sawtooth < x"dff" then   pst_out <= x"8c";
      elsif sawtooth < x"e00" then   pst_out <= x"9f";
      elsif sawtooth < x"e3e" then   pst_out <= x"00";
      elsif sawtooth < x"e40" then   pst_out <= x"80";
      elsif sawtooth < x"e5e" then   pst_out <= x"00";
      elsif sawtooth < x"e60" then   pst_out <= x"80";
      elsif sawtooth < x"e66" then   pst_out <= x"00";
      elsif sawtooth < x"e67" then   pst_out <= x"80";
      elsif sawtooth < x"e6a" then   pst_out <= x"00";
      elsif sawtooth < x"e80" then   pst_out <= x"80";
      elsif sawtooth < x"e82" then   pst_out <= x"00";
      elsif sawtooth < x"e83" then   pst_out <= x"80";
      elsif sawtooth < x"e85" then   pst_out <= x"00";
      elsif sawtooth < x"e89" then   pst_out <= x"80";
      elsif sawtooth < x"e8a" then   pst_out <= x"00";
      elsif sawtooth < x"eee" then   pst_out <= x"80";
      elsif sawtooth < x"eff" then   pst_out <= x"c0";
      elsif sawtooth < x"f00" then   pst_out <= x"cf";
      elsif sawtooth < x"f6f" then   pst_out <= x"c0";
      elsif sawtooth < x"f70" then   pst_out <= x"e0";
      elsif sawtooth < x"f74" then   pst_out <= x"c0";
      elsif sawtooth < x"f7f" then   pst_out <= x"e0";
      elsif sawtooth < x"f80" then   pst_out <= x"e3";
      elsif sawtooth < x"fb6" then   pst_out <= x"e0";
      elsif sawtooth < x"fda" then   pst_out <= x"f0";
      elsif sawtooth < x"feb" then   pst_out <= x"f8";
      elsif sawtooth < x"ff5" then   pst_out <= x"fc";
      elsif sawtooth < x"ff9" then   pst_out <= x"fe";
      else  pst_out <= x"ff";
      end if;
      
      
    end if;
  end process;
  
end sequential;
