module UART_TX_CTRL (input CLK, input SEND, output READY, output UART_TX, input [7:0] DATA, input [15:0] BIT_TMR_MAX);
   

endmodule
