library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

--
entity kickstart is
  port (Clk : in std_logic;
        address : in std_logic_vector(13 downto 0);
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        we : in std_logic;
        -- chip select, active low       
        cs : in std_logic;
        data_i : in std_logic_vector(7 downto 0);
        data_o : out std_logic_vector(7 downto 0)
        );
end kickstart;

architecture Behavioral of kickstart is

-- 16K x 8bit pre-initialised RAM
  type ram_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal ram : ram_t := (x"78",x"D8",x"03",x"A9",x"00",x"8D",x"17",x"D0",x"A9",x"00",x"5B",x"A0",x"01",x"2B",x"A2",x"FF",x"9A",x"A9",x"7F",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"A9",x"00",x"8D",x"1A",x"D0",x"4C",x"21",x"80",x"A9",x"7F",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"A9",x"00",x"8D",x"19",x"D0",x"38",x"20",x"1E",x"8C",x"20",x"78",x"89",x"20",x"8A",x"8A",x"20",x"A3",x"89",x"A2",x"FB",x"A0",x"8C",x"20",x"EA",x"8A",x"EE",x"01",x"CF",x"20",x"31",x"8C",x"AD",x"F1",x"D6",x"29",x"02",x"F0",x"06",x"20",x"90",x"8C",x"4C",x"4F",x"80",x"A2",x"73",x"A0",x"8D",x"20",x"EA",x"8A",x"20",x"10",x"87",x"B0",x"03",x"4C",x"5C",x"80",x"A2",x"13",x"A0",x"8E",x"20",x"EA",x"8A",x"A9",x"3E",x"8D",x"C0",x"07",x"20",x"B7",x"87",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"53",x"04",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"4B",x"04",x"A2",x"3B",x"A0",x"8E",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"C2",x"DF",x"20",x"32",x"8B",x"AB",x"C9",x"DF",x"9C",x"0B",x"CF",x"20",x"32",x"8B",x"AB",x"C8",x"DF",x"9C",x"0A",x"CF",x"20",x"32",x"8B",x"AB",x"C7",x"DF",x"9C",x"09",x"CF",x"20",x"32",x"8B",x"AB",x"C6",x"DF",x"9C",x"08",x"CF",x"20",x"32",x"8B",x"AB",x"CD",x"DF",x"20",x"32",x"8B",x"AB",x"CC",x"DF",x"20",x"32",x"8B",x"AB",x"CB",x"DF",x"20",x"32",x"8B",x"AB",x"CA",x"DF",x"20",x"32",x"8B",x"A2",x"03",x"BD",x"08",x"CF",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"20",x"81",x"88",x"20",x"C5",x"87",x"93",x"DF",x"03",x"A9",x"3E",x"8D",x"C1",x"07",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"DF",x"03",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"D7",x"03",x"A2",x"63",x"A0",x"8E",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"0D",x"DE",x"20",x"32",x"8B",x"AB",x"0F",x"DE",x"20",x"32",x"8B",x"AB",x"0E",x"DE",x"20",x"32",x"8B",x"AB",x"2F",x"DE",x"20",x"32",x"8B",x"AB",x"2E",x"DE",x"20",x"32",x"8B",x"AB",x"2D",x"DE",x"20",x"32",x"8B",x"AB",x"2C",x"DE",x"20",x"32",x"8B",x"AD",x"11",x"DE",x"D3",x"9E",x"03",x"A2",x"03",x"BD",x"0E",x"DE",x"9D",x"10",x"CF",x"9D",x"0C",x"CF",x"BD",x"2C",x"DE",x"9D",x"14",x"CF",x"CA",x"10",x"EE",x"A9",x"00",x"8D",x"12",x"CF",x"8D",x"13",x"CF",x"8D",x"0E",x"CF",x"8D",x"0F",x"CF",x"AC",x"10",x"DE",x"F0",x"18",x"A2",x"00",x"18",x"08",x"28",x"BD",x"10",x"CF",x"7D",x"24",x"DE",x"9D",x"10",x"CF",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"88",x"D0",x"E8",x"38",x"A2",x"03",x"BD",x"20",x"DE",x"FD",x"10",x"CF",x"9D",x"1C",x"CF",x"9D",x"20",x"CF",x"CA",x"10",x"F1",x"AD",x"0D",x"DE",x"8D",x"24",x"CF",x"A8",x"29",x"FE",x"F0",x"14",x"A2",x"03",x"18",x"BD",x"20",x"CF",x"6A",x"9D",x"20",x"CF",x"CA",x"10",x"F6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"AD",x"23",x"CF",x"0D",x"22",x"CF",x"F3",x"25",x"03",x"A2",x"8B",x"A0",x"8E",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"13",x"CF",x"20",x"32",x"8B",x"AB",x"12",x"CF",x"20",x"32",x"8B",x"AB",x"11",x"CF",x"20",x"32",x"8B",x"AB",x"10",x"CF",x"20",x"32",x"8B",x"AB",x"1F",x"CF",x"20",x"32",x"8B",x"AB",x"1E",x"CF",x"20",x"32",x"8B",x"AB",x"1D",x"CF",x"20",x"32",x"8B",x"AB",x"1C",x"CF",x"20",x"32",x"8B",x"AB",x"23",x"CF",x"20",x"32",x"8B",x"AB",x"22",x"CF",x"20",x"32",x"8B",x"AB",x"21",x"CF",x"20",x"32",x"8B",x"AB",x"20",x"CF",x"20",x"32",x"8B",x"A2",x"03",x"BD",x"2C",x"DE",x"9D",x"18",x"CF",x"9D",x"4A",x"CF",x"CA",x"10",x"F4",x"20",x"E5",x"84",x"20",x"F4",x"84",x"93",x"B0",x"02",x"20",x"09",x"85",x"93",x"75",x"00",x"A2",x"00",x"BD",x"29",x"CF",x"20",x"DA",x"84",x"DD",x"99",x"91",x"D0",x"ED",x"E8",x"E0",x"0B",x"D0",x"F0",x"A2",x"0B",x"A0",x"91",x"20",x"EA",x"8A",x"A9",x"00",x"85",x"FB",x"85",x"FD",x"85",x"FE",x"A9",x"40",x"85",x"FC",x"20",x"58",x"85",x"20",x"78",x"86",x"20",x"72",x"85",x"90",x"44",x"A3",x"00",x"B9",x"00",x"DE",x"EA",x"92",x"FB",x"1B",x"D0",x"F7",x"E3",x"FC",x"B9",x"00",x"DF",x"EA",x"92",x"FB",x"1B",x"D0",x"F7",x"E3",x"FC",x"20",x"83",x"85",x"B0",x"E3",x"A2",x"5B",x"A0",x"91",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"FE",x"00",x"20",x"32",x"8B",x"AB",x"FD",x"00",x"20",x"32",x"8B",x"AB",x"FC",x"00",x"20",x"32",x"8B",x"AB",x"FB",x"00",x"20",x"32",x"8B",x"20",x"00",x"40",x"4C",x"92",x"82",x"A2",x"33",x"A0",x"91",x"20",x"EA",x"8A",x"A9",x"3E",x"8D",x"C2",x"07",x"A9",x"00",x"8D",x"8B",x"D6",x"20",x"E5",x"84",x"20",x"F4",x"84",x"93",x"1C",x"02",x"20",x"09",x"85",x"93",x"E6",x"00",x"A2",x"00",x"BD",x"29",x"CF",x"20",x"DA",x"84",x"DD",x"8E",x"91",x"D0",x"ED",x"E8",x"E0",x"0B",x"D0",x"F0",x"A2",x"1B",x"A0",x"90",x"20",x"EA",x"8A",x"20",x"58",x"85",x"20",x"78",x"86",x"20",x"81",x"88",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"8C",x"D6",x"CA",x"10",x"F7",x"20",x"58",x"85",x"A2",x"03",x"BD",x"4A",x"CF",x"9D",x"4F",x"CF",x"CA",x"10",x"F7",x"A9",x"00",x"8D",x"55",x"CF",x"8D",x"56",x"CF",x"A9",x"40",x"8D",x"53",x"CF",x"A9",x"06",x"8D",x"54",x"CF",x"AB",x"24",x"CF",x"6B",x"29",x"01",x"D0",x"0C",x"6B",x"4A",x"4B",x"4E",x"54",x"CF",x"6E",x"53",x"CF",x"4C",x"FB",x"82",x"A2",x"03",x"BD",x"4F",x"CF",x"DD",x"4A",x"CF",x"D0",x"5A",x"CA",x"10",x"F5",x"EE",x"55",x"CF",x"D0",x"03",x"EE",x"56",x"CF",x"18",x"AD",x"4F",x"CF",x"69",x"01",x"8D",x"4F",x"CF",x"AD",x"50",x"CF",x"69",x"00",x"8D",x"50",x"CF",x"AD",x"51",x"CF",x"69",x"00",x"8D",x"51",x"CF",x"AD",x"52",x"CF",x"69",x"00",x"8D",x"52",x"CF",x"20",x"C2",x"85",x"B0",x"C5",x"AD",x"53",x"CF",x"CD",x"55",x"CF",x"D0",x"17",x"AD",x"54",x"CF",x"CD",x"56",x"CF",x"D0",x"0F",x"A9",x"07",x"8D",x"8B",x"D6",x"A2",x"93",x"A0",x"90",x"20",x"EA",x"8A",x"4C",x"97",x"83",x"A2",x"43",x"A0",x"90",x"20",x"EA",x"8A",x"4C",x"97",x"83",x"EE",x"20",x"D0",x"A2",x"00",x"BD",x"4F",x"CF",x"9D",x"28",x"04",x"BD",x"4A",x"CF",x"9D",x"30",x"04",x"E8",x"E0",x"04",x"D0",x"EF",x"A2",x"6B",x"A0",x"90",x"20",x"EA",x"8A",x"4C",x"97",x"83",x"A2",x"F3",x"A0",x"8F",x"20",x"EA",x"8A",x"20",x"B6",x"88",x"90",x"0A",x"A2",x"23",x"A0",x"8D",x"20",x"EA",x"8A",x"4C",x"57",x"8B",x"A2",x"4B",x"A0",x"8D",x"20",x"EA",x"8A",x"20",x"E5",x"84",x"20",x"F4",x"84",x"93",x"0B",x"01",x"20",x"09",x"85",x"B0",x"21",x"A2",x"0B",x"BD",x"83",x"91",x"9D",x"F6",x"90",x"CA",x"D0",x"F7",x"A2",x"E3",x"A0",x"90",x"20",x"EA",x"8A",x"20",x"6E",x"87",x"20",x"6E",x"87",x"20",x"6E",x"87",x"20",x"6E",x"87",x"4C",x"C0",x"84",x"A2",x"00",x"BD",x"29",x"CF",x"20",x"DA",x"84",x"DD",x"83",x"91",x"D0",x"CD",x"E8",x"E0",x"0B",x"D0",x"F0",x"20",x"58",x"85",x"A9",x"3E",x"8D",x"C3",x"07",x"A2",x"DB",x"A0",x"8E",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"4D",x"CF",x"20",x"32",x"8B",x"AB",x"4C",x"CF",x"20",x"32",x"8B",x"AB",x"4B",x"CF",x"20",x"32",x"8B",x"AB",x"4A",x"CF",x"20",x"32",x"8B",x"20",x"72",x"85",x"93",x"9D",x"00",x"A2",x"2B",x"A0",x"8F",x"20",x"EA",x"8A",x"A9",x"00",x"8D",x"06",x"CF",x"8D",x"07",x"CF",x"A9",x"80",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"AD",x"06",x"CF",x"0A",x"85",x"FB",x"AD",x"06",x"CF",x"4A",x"4A",x"4A",x"4A",x"4A",x"4A",x"4A",x"85",x"FC",x"A5",x"FB",x"18",x"69",x"C0",x"85",x"FB",x"A5",x"FC",x"69",x"01",x"09",x"40",x"AA",x"A5",x"FB",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A2",x"00",x"BD",x"00",x"DE",x"9D",x"00",x"40",x"BD",x"00",x"DF",x"9D",x"00",x"41",x"E8",x"D0",x"F1",x"A9",x"00",x"AA",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A9",x"00",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"EE",x"06",x"CF",x"D0",x"03",x"EE",x"07",x"CF",x"AD",x"07",x"CF",x"C9",x"02",x"F0",x"21",x"EE",x"20",x"D0",x"20",x"83",x"85",x"B0",x"93",x"AD",x"06",x"CF",x"D0",x"14",x"AD",x"07",x"CF",x"C9",x"01",x"D0",x"0D",x"20",x"E9",x"88",x"A2",x"23",x"A0",x"8D",x"20",x"EA",x"8A",x"4C",x"57",x"8B",x"A2",x"53",x"A0",x"8F",x"20",x"EA",x"8A",x"A2",x"03",x"A0",x"8F",x"20",x"EA",x"8A",x"A2",x"C3",x"A0",x"8D",x"20",x"EA",x"8A",x"20",x"6E",x"87",x"4C",x"00",x"80",x"A2",x"EB",x"A0",x"8D",x"20",x"EA",x"8A",x"20",x"6E",x"87",x"4C",x"00",x"80",x"C9",x"60",x"90",x"06",x"C9",x"7A",x"B0",x"02",x"29",x"5F",x"60",x"A2",x"00",x"BD",x"18",x"CF",x"9D",x"25",x"CF",x"E8",x"E0",x"04",x"D0",x"F5",x"38",x"60",x"A2",x"00",x"BD",x"25",x"CF",x"9D",x"4A",x"CF",x"E8",x"E0",x"04",x"D0",x"F5",x"A9",x"00",x"8D",x"49",x"CF",x"4C",x"72",x"85",x"AD",x"49",x"CF",x"C9",x"10",x"90",x"0B",x"A9",x"00",x"8D",x"49",x"CF",x"20",x"83",x"85",x"B0",x"01",x"60",x"A0",x"00",x"AD",x"49",x"CF",x"29",x"08",x"D0",x"1A",x"AD",x"49",x"CF",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DE",x"99",x"29",x"CF",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CF",x"38",x"60",x"AD",x"49",x"CF",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DF",x"99",x"29",x"CF",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CF",x"38",x"60",x"AD",x"3D",x"CF",x"8D",x"4C",x"CF",x"AD",x"3E",x"CF",x"8D",x"4D",x"CF",x"AD",x"43",x"CF",x"8D",x"4A",x"CF",x"AD",x"44",x"CF",x"8D",x"4B",x"CF",x"38",x"60",x"A9",x"00",x"8D",x"4E",x"CF",x"20",x"78",x"86",x"B0",x"01",x"60",x"20",x"81",x"88",x"4C",x"C5",x"87",x"20",x"4D",x"88",x"EE",x"4E",x"CF",x"AD",x"4E",x"CF",x"CD",x"24",x"CF",x"D0",x"20",x"A9",x"00",x"8D",x"4E",x"CF",x"20",x"C2",x"85",x"B0",x"01",x"60",x"20",x"78",x"86",x"20",x"81",x"88",x"08",x"AD",x"F1",x"D6",x"29",x"10",x"F0",x"06",x"20",x"EA",x"86",x"20",x"6E",x"87",x"28",x"4C",x"C5",x"87",x"49",x"54",x"53",x"20",x"52",x"49",x"47",x"48",x"54",x"20",x"48",x"45",x"52",x"45",x"A2",x"00",x"BD",x"4A",x"CF",x"9D",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F5",x"A0",x"07",x"18",x"6E",x"84",x"D6",x"6E",x"83",x"D6",x"6E",x"82",x"D6",x"6E",x"81",x"D6",x"88",x"D0",x"F0",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"0C",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"20",x"81",x"88",x"20",x"C5",x"87",x"90",x"63",x"AD",x"4A",x"CF",x"0A",x"0A",x"AA",x"A0",x"00",x"AD",x"4A",x"CF",x"29",x"40",x"D0",x"0E",x"BD",x"00",x"DE",x"99",x"4A",x"CF",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"80",x"0C",x"BD",x"00",x"DF",x"99",x"4A",x"CF",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"AD",x"4D",x"CF",x"29",x"0F",x"8D",x"4D",x"CF",x"AD",x"4D",x"CF",x"0D",x"4C",x"CF",x"0D",x"4B",x"CF",x"0D",x"4A",x"CF",x"C9",x"00",x"F0",x"22",x"AD",x"4D",x"CF",x"C9",x"0F",x"D0",x"19",x"AD",x"4C",x"CF",x"C9",x"FF",x"D0",x"12",x"AD",x"4B",x"CF",x"C9",x"FF",x"D0",x"0B",x"AD",x"4A",x"CF",x"C9",x"FF",x"F0",x"06",x"C9",x"F7",x"F0",x"02",x"38",x"60",x"18",x"60",x"A2",x"03",x"BD",x"4A",x"CF",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A2",x"00",x"38",x"08",x"28",x"BD",x"81",x"D6",x"FD",x"14",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"AD",x"24",x"CF",x"A8",x"29",x"FE",x"F0",x"14",x"18",x"2E",x"81",x"D6",x"2E",x"82",x"D6",x"2E",x"83",x"D6",x"2E",x"84",x"D6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"A2",x"00",x"BD",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"10",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"38",x"60",x"A2",x"B3",x"A0",x"8E",x"20",x"EA",x"8A",x"A0",x"00",x"A2",x"03",x"BD",x"4A",x"CF",x"4B",x"DA",x"20",x"32",x"8B",x"FA",x"CA",x"10",x"F4",x"A2",x"03",x"BD",x"81",x"D6",x"4B",x"DA",x"20",x"32",x"8B",x"FA",x"CA",x"10",x"F4",x"60",x"20",x"2E",x"87",x"B0",x"01",x"60",x"A2",x"9B",x"A0",x"8D",x"20",x"EA",x"8A",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"4C",x"C5",x"87",x"A9",x"42",x"8D",x"80",x"D6",x"A9",x"00",x"8D",x"80",x"D6",x"20",x"8D",x"87",x"20",x"9B",x"87",x"B0",x"03",x"D0",x"F9",x"60",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"8D",x"87",x"20",x"9B",x"87",x"B0",x"03",x"D0",x"F9",x"60",x"20",x"6E",x"87",x"20",x"B7",x"87",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"8D",x"87",x"AD",x"80",x"D6",x"20",x"9B",x"87",x"B0",x"03",x"D0",x"F6",x"60",x"38",x"60",x"20",x"8D",x"87",x"20",x"90",x"8C",x"EE",x"20",x"D0",x"20",x"C1",x"8C",x"CE",x"20",x"D0",x"EE",x"00",x"03",x"D0",x"F2",x"EE",x"01",x"03",x"D0",x"ED",x"EE",x"02",x"03",x"D0",x"E8",x"60",x"A9",x"00",x"8D",x"00",x"03",x"8D",x"01",x"03",x"A9",x"F7",x"8D",x"02",x"03",x"60",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"13",x"EE",x"00",x"03",x"D0",x"0C",x"EE",x"01",x"03",x"D0",x"07",x"EE",x"02",x"03",x"D0",x"02",x"A9",x"00",x"18",x"60",x"38",x"60",x"A9",x"81",x"8D",x"80",x"D6",x"38",x"60",x"A9",x"82",x"8D",x"80",x"D6",x"38",x"60",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"3D",x"4C",x"DE",x"87",x"A2",x"F0",x"A0",x"00",x"A3",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"E8",x"D0",x"F7",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"8D",x"87",x"20",x"9B",x"87",x"B0",x"05",x"D0",x"F9",x"4C",x"03",x"88",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"EF",x"AD",x"88",x"D6",x"AD",x"89",x"D6",x"C9",x"02",x"D0",x"CE",x"38",x"60",x"20",x"2E",x"87",x"4C",x"DE",x"87",x"18",x"60",x"A2",x"7B",x"A0",x"8F",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"4D",x"CF",x"20",x"32",x"8B",x"AB",x"4C",x"CF",x"20",x"32",x"8B",x"AB",x"4B",x"CF",x"20",x"32",x"8B",x"AB",x"4A",x"CF",x"4C",x"32",x"8B",x"A2",x"A3",x"A0",x"8F",x"20",x"EA",x"8A",x"A0",x"00",x"AB",x"84",x"D6",x"20",x"32",x"8B",x"AB",x"83",x"D6",x"20",x"32",x"8B",x"AB",x"82",x"D6",x"20",x"32",x"8B",x"AB",x"81",x"D6",x"4C",x"32",x"8B",x"AD",x"80",x"D6",x"29",x"10",x"D0",x"1A",x"AD",x"82",x"D6",x"18",x"69",x"02",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"69",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"69",x"00",x"8D",x"84",x"D6",x"60",x"EE",x"81",x"D6",x"90",x"0D",x"EE",x"82",x"D6",x"90",x"08",x"EE",x"83",x"D6",x"90",x"03",x"EE",x"84",x"D6",x"60",x"AD",x"80",x"D6",x"29",x"10",x"F0",x"01",x"60",x"AD",x"83",x"D6",x"8D",x"84",x"D6",x"AD",x"82",x"D6",x"8D",x"83",x"D6",x"AD",x"81",x"D6",x"8D",x"82",x"D6",x"A9",x"00",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"0A",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"2A",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"2A",x"8D",x"84",x"D6",x"60",x"AD",x"F1",x"D6",x"29",x"20",x"D0",x"2A",x"AD",x"88",x"91",x"C9",x"20",x"D0",x"23",x"20",x"13",x"89",x"20",x"FF",x"88",x"AD",x"00",x"40",x"CD",x"02",x"CF",x"D0",x"15",x"AD",x"01",x"40",x"CD",x"03",x"CF",x"D0",x"0D",x"AD",x"02",x"40",x"CD",x"04",x"CF",x"D0",x"05",x"20",x"0D",x"8C",x"38",x"60",x"18",x"60",x"20",x"FF",x"88",x"AD",x"02",x"CF",x"8D",x"00",x"40",x"AD",x"03",x"CF",x"8D",x"01",x"40",x"AD",x"04",x"CF",x"8D",x"02",x"40",x"60",x"A9",x"80",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"A9",x"C0",x"A2",x"CF",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"60",x"A9",x"03",x"8D",x"02",x"CF",x"8D",x"03",x"CF",x"8D",x"04",x"CF",x"8D",x"05",x"CF",x"A9",x"08",x"8D",x"00",x"CF",x"AD",x"00",x"CF",x"38",x"E9",x"01",x"4A",x"4A",x"09",x"C0",x"AA",x"AD",x"00",x"CF",x"38",x"E9",x"01",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A9",x"00",x"85",x"FB",x"A9",x"40",x"85",x"FC",x"A0",x"00",x"AD",x"02",x"CF",x"18",x"71",x"FB",x"8D",x"02",x"CF",x"90",x"08",x"EE",x"03",x"CF",x"90",x"03",x"EE",x"04",x"CF",x"C8",x"D0",x"EA",x"E6",x"FC",x"A5",x"FC",x"C9",x"80",x"D0",x"E0",x"EE",x"00",x"CF",x"AD",x"00",x"CF",x"C9",x"10",x"D0",x"B1",x"4C",x"0D",x"8C",x"A9",x"40",x"8D",x"30",x"D0",x"A9",x"00",x"8D",x"31",x"D0",x"8D",x"20",x"D0",x"8D",x"21",x"D0",x"8D",x"54",x"D0",x"A9",x"14",x"8D",x"18",x"D0",x"A9",x"1B",x"8D",x"11",x"D0",x"A9",x"C8",x"8D",x"16",x"D0",x"A9",x"FF",x"8D",x"01",x"DD",x"8D",x"00",x"DD",x"60",x"A9",x"04",x"8D",x"30",x"D0",x"A9",x"FF",x"8D",x"70",x"D0",x"A9",x"00",x"8D",x"00",x"D1",x"8D",x"00",x"D2",x"8D",x"00",x"D3",x"A9",x"FF",x"8D",x"01",x"D1",x"8D",x"01",x"D2",x"8D",x"01",x"D3",x"A9",x"BA",x"8D",x"02",x"D1",x"A9",x"13",x"8D",x"02",x"D2",x"A9",x"62",x"8D",x"02",x"D3",x"A9",x"66",x"8D",x"03",x"D1",x"A9",x"AD",x"8D",x"03",x"D2",x"A9",x"FF",x"8D",x"03",x"D3",x"A9",x"BB",x"8D",x"04",x"D1",x"A9",x"F3",x"8D",x"04",x"D2",x"A9",x"8B",x"8D",x"04",x"D3",x"A9",x"55",x"8D",x"05",x"D1",x"A9",x"EC",x"8D",x"05",x"D2",x"A9",x"85",x"8D",x"05",x"D3",x"A9",x"D1",x"8D",x"06",x"D1",x"A9",x"E0",x"8D",x"06",x"D2",x"A9",x"79",x"8D",x"06",x"D3",x"A9",x"AE",x"8D",x"07",x"D1",x"A9",x"5F",x"8D",x"07",x"D2",x"A9",x"C7",x"8D",x"07",x"D3",x"A9",x"9B",x"8D",x"08",x"D1",x"A9",x"47",x"8D",x"08",x"D2",x"A9",x"81",x"8D",x"08",x"D3",x"A9",x"87",x"8D",x"09",x"D1",x"A9",x"37",x"8D",x"09",x"D2",x"A9",x"00",x"8D",x"09",x"D3",x"A9",x"DD",x"8D",x"0A",x"D1",x"A9",x"39",x"8D",x"0A",x"D2",x"A9",x"78",x"8D",x"0A",x"D3",x"A9",x"B5",x"8D",x"0B",x"D1",x"8D",x"0B",x"D2",x"8D",x"0B",x"D3",x"A9",x"B8",x"8D",x"0C",x"D1",x"8D",x"0C",x"D2",x"8D",x"0C",x"D3",x"A9",x"0B",x"8D",x"0D",x"D1",x"A9",x"4F",x"8D",x"0D",x"D2",x"A9",x"CA",x"8D",x"0D",x"D3",x"A9",x"AA",x"8D",x"0E",x"D1",x"A9",x"D9",x"8D",x"0E",x"D2",x"A9",x"FE",x"8D",x"0E",x"D3",x"A9",x"8B",x"8D",x"0F",x"D1",x"8D",x"0F",x"D2",x"8D",x"0F",x"D3",x"60",x"A9",x"01",x"0C",x"30",x"D0",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"8D",x"05",x"D7",x"A9",x"00",x"8D",x"06",x"D7",x"A9",x"8A",x"8D",x"01",x"D7",x"A9",x"BB",x"8D",x"00",x"D7",x"A9",x"00",x"8D",x"05",x"D7",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"00",x"8D",x"01",x"CF",x"60",x"07",x"E8",x"03",x"20",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"07",x"D0",x"07",x"01",x"00",x"00",x"00",x"D8",x"80",x"00",x"00",x"00",x"00",x"10",x"A4",x"91",x"0F",x"00",x"C0",x"00",x"00",x"00",x"48",x"A2",x"CB",x"A0",x"8F",x"20",x"EA",x"8A",x"A0",x"00",x"FB",x"4C",x"32",x"8B",x"86",x"FB",x"84",x"FC",x"A9",x"00",x"85",x"FD",x"A9",x"04",x"85",x"FE",x"AE",x"01",x"CF",x"E0",x"00",x"F0",x"22",x"18",x"A5",x"FD",x"69",x"28",x"85",x"FD",x"A5",x"FE",x"69",x"00",x"85",x"FE",x"C9",x"07",x"90",x"0E",x"A5",x"FD",x"C9",x"E8",x"90",x"08",x"A9",x"00",x"85",x"FD",x"A9",x"04",x"85",x"FE",x"CA",x"D0",x"DA",x"A0",x"27",x"B1",x"FB",x"C9",x"40",x"90",x"02",x"29",x"1F",x"91",x"FD",x"88",x"10",x"F3",x"EE",x"01",x"CF",x"60",x"6B",x"4A",x"4A",x"4A",x"4A",x"20",x"3D",x"8B",x"6B",x"29",x"0F",x"AA",x"B1",x"FD",x"C9",x"24",x"F0",x"06",x"C8",x"C0",x"28",x"D0",x"F5",x"60",x"8A",x"09",x"30",x"C9",x"3A",x"90",x"02",x"E9",x"39",x"91",x"FD",x"C8",x"60",x"AD",x"F1",x"D6",x"10",x"0C",x"A2",x"BB",x"A0",x"90",x"20",x"EA",x"8A",x"AD",x"F1",x"D6",x"30",x"FB",x"A9",x"82",x"8D",x"80",x"D6",x"A2",x"00",x"8A",x"9D",x"00",x"08",x"E8",x"D0",x"FA",x"A9",x"00",x"8D",x"40",x"D6",x"8D",x"41",x"D6",x"8D",x"42",x"D6",x"8D",x"43",x"D6",x"8D",x"44",x"D6",x"A9",x"FF",x"8D",x"45",x"D6",x"A9",x"01",x"8D",x"46",x"D6",x"A9",x"F7",x"8D",x"47",x"D6",x"A2",x"FC",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"DC",x"8B",x"AD",x"00",x"BC",x"8D",x"48",x"D6",x"A2",x"FD",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"DC",x"8B",x"AD",x"00",x"BC",x"8D",x"49",x"D6",x"A9",x"00",x"8D",x"4A",x"D6",x"8D",x"4B",x"D6",x"8D",x"4C",x"D6",x"8D",x"4D",x"D6",x"8D",x"4E",x"D6",x"8D",x"4F",x"D6",x"A9",x"3F",x"8D",x"50",x"D6",x"8D",x"51",x"D6",x"A9",x"00",x"8D",x"52",x"D6",x"8D",x"7F",x"D6",x"8D",x"05",x"D7",x"A9",x"FF",x"8D",x"06",x"D7",x"8E",x"05",x"8C",x"8C",x"06",x"8C",x"9C",x"07",x"8C",x"A9",x"8C",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"02",x"8D",x"00",x"D7",x"60",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"BC",x"0F",x"00",x"00",x"A9",x"00",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"AA",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"60",x"B0",x"06",x"A9",x"00",x"8D",x"2F",x"D0",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"60",x"A9",x"FF",x"8D",x"03",x"DC",x"A9",x"00",x"8D",x"02",x"DC",x"A9",x"FE",x"8D",x"01",x"DC",x"A9",x"20",x"AE",x"00",x"DC",x"E0",x"7F",x"D0",x"02",x"A9",x"31",x"E0",x"EF",x"D0",x"02",x"A9",x"39",x"E0",x"F7",x"D0",x"02",x"A9",x"37",x"E0",x"FB",x"D0",x"02",x"A9",x"35",x"E0",x"FD",x"D0",x"02",x"A9",x"33",x"A2",x"F7",x"8E",x"01",x"DC",x"AE",x"00",x"DC",x"E0",x"7F",x"D0",x"02",x"A9",x"32",x"E0",x"EF",x"D0",x"02",x"A9",x"30",x"E0",x"F7",x"D0",x"02",x"A9",x"38",x"E0",x"FB",x"D0",x"02",x"A9",x"36",x"E0",x"FD",x"D0",x"02",x"A9",x"34",x"8D",x"88",x"91",x"8D",x"27",x"04",x"60",x"AD",x"F1",x"D6",x"29",x"01",x"D0",x"01",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"A9",x"FF",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A9",x"80",x"A2",x"8D",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"AD",x"E1",x"D6",x"4A",x"29",x"02",x"09",x"01",x"8D",x"E1",x"D6",x"AD",x"E1",x"D6",x"29",x"20",x"D0",x"01",x"60",x"AD",x"E1",x"D6",x"29",x"04",x"4A",x"09",x"01",x"8D",x"E1",x"D6",x"AD",x"10",x"68",x"C9",x"45",x"D0",x"1F",x"AD",x"19",x"68",x"C9",x"11",x"D0",x"18",x"AD",x"26",x"68",x"C9",x"11",x"D0",x"11",x"AD",x"27",x"68",x"C9",x"9F",x"D0",x"0A",x"AD",x"2C",x"68",x"C9",x"A9",x"D0",x"03",x"20",x"2C",x"68",x"60",x"43",x"36",x"35",x"47",x"53",x"20",x"4B",x"49",x"43",x"4B",x"53",x"54",x"41",x"52",x"54",x"20",x"56",x"30",x"30",x"2E",x"30",x"30",x"20",x"50",x"52",x"45",x"2D",x"41",x"4C",x"50",x"48",x"41",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"4F",x"4D",x"20",x"43",x"48",x"45",x"43",x"4B",x"53",x"55",x"4D",x"20",x"4F",x"4B",x"20",x"2D",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"4F",x"4D",x"20",x"43",x"48",x"45",x"43",x"4B",x"53",x"55",x"4D",x"20",x"46",x"41",x"49",x"4C",x"20",x"2D",x"20",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"52",x"4F",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"2E",x"2E",x"2E",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"46",x"4F",x"55",x"4E",x"44",x"20",x"41",x"4E",x"44",x"20",x"52",x"45",x"53",x"45",x"54",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"20",x"43",x"41",x"52",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"44",x"20",x"4D",x"42",x"52",x"20",x"4F",x"52",x"20",x"44",x"4F",x"53",x"20",x"42",x"4F",x"4F",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"2E",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"45",x"41",x"44",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"54",x"41",x"42",x"4C",x"45",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"31",x"28",x"24",x"24",x"29",x"20",x"40",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"2C",x"20",x"53",x"49",x"5A",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"46",x"53",x"20",x"53",x"50",x"43",x"3A",x"24",x"24",x"20",x"52",x"53",x"56",x"53",x"45",x"43",x"3A",x"24",x"24",x"24",x"24",x"20",x"52",x"53",x"56",x"43",x"4C",x"55",x"53",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"53",x"59",x"53",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"44",x"41",x"54",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"43",x"4C",x"55",x"53",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"2D",x"3E",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"3A",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"46",x"4F",x"55",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"20",x"3D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4F",x"50",x"45",x"4E",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"20",x"46",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"20",x"20",x"20",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"2E",x"2E",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"20",x"57",x"52",x"4F",x"4E",x"47",x"20",x"53",x"49",x"5A",x"45",x"3A",x"20",x"4D",x"55",x"53",x"54",x"20",x"42",x"45",x"20",x"31",x"32",x"38",x"4B",x"42",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"58",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"3D",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"58",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"3D",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"48",x"45",x"43",x"4B",x"50",x"4F",x"49",x"4E",x"54",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"43",x"41",x"4E",x"4E",x"4F",x"54",x"20",x"46",x"49",x"4E",x"44",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"2D",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"20",x"44",x"49",x"53",x"4B",x"4C",x"45",x"53",x"53",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"40",x"20",x"49",x"4E",x"54",x"45",x"52",x"4E",x"41",x"4C",x"20",x"46",x"30",x"31",x"31",x"20",x"44",x"52",x"49",x"56",x"45",x"46",x"41",x"49",x"4C",x"3A",x"20",x"43",x"36",x"34",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"49",x"53",x"20",x"4E",x"4F",x"54",x"20",x"38",x"31",x"39",x"32",x"30",x"30",x"20",x"42",x"59",x"54",x"45",x"53",x"20",x"4C",x"4F",x"4E",x"47",x"46",x"41",x"49",x"4C",x"3A",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"49",x"53",x"20",x"46",x"52",x"41",x"47",x"4D",x"45",x"4E",x"54",x"45",x"44",x"3A",x"20",x"44",x"45",x"46",x"52",x"41",x"47",x"20",x"49",x"54",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"53",x"55",x"43",x"43",x"45",x"53",x"53",x"46",x"55",x"4C",x"4C",x"59",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"45",x"4C",x"45",x"41",x"53",x"45",x"20",x"53",x"57",x"31",x"35",x"20",x"54",x"4F",x"20",x"43",x"4F",x"4E",x"54",x"49",x"4E",x"55",x"45",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"2E",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"46",x"49",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"43",x"36",x"35",x"47",x"53",x"58",x"58",x"58",x"52",x"4F",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"4B",x"49",x"43",x"4B",x"55",x"50",x"2E",x"47",x"36",x"35",x"20",x"49",x"4E",x"54",x"4F",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"4F",x"20",x"4B",x"49",x"43",x"4B",x"55",x"50",x"2E",x"47",x"36",x"35",x"20",x"54",x"4F",x"20",x"4C",x"4F",x"41",x"44",x"20",x"28",x"4F",x"52",x"20",x"42",x"52",x"4F",x"4B",x"45",x"4E",x"29",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4B",x"49",x"43",x"4B",x"55",x"50",x"20",x"4C",x"4F",x"41",x"44",x"45",x"44",x"20",x"54",x"4F",x"20",x"30",x"30",x"30",x"30",x"34",x"30",x"30",x"30",x"20",x"2D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"43",x"36",x"35",x"47",x"53",x"20",x"20",x"20",x"52",x"4F",x"4D",x"43",x"36",x"35",x"47",x"53",x"20",x"20",x"20",x"44",x"38",x"31",x"4B",x"49",x"43",x"4B",x"55",x"50",x"20",x"20",x"47",x"36",x"35",x"BA",x"8E",x"5A",x"CF",x"A9",x"93",x"20",x"D2",x"FF",x"38",x"20",x"DC",x"C6",x"78",x"20",x"AC",x"C6",x"4F",x"50",x"45",x"4E",x"49",x"4E",x"47",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"2E",x"2E",x"2E",x"0D",x"00",x"20",x"5E",x"C5",x"B0",x"03",x"4C",x"24",x"C0",x"20",x"AC",x"C6",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"54",x"41",x"42",x"4C",x"45",x"2E",x"2E",x"2E",x"0D",x"00",x"20",x"EC",x"C5",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"DB",x"02",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"D3",x"02",x"A0",x"00",x"AB",x"C9",x"DF",x"9C",x"0B",x"CF",x"AB",x"C8",x"DF",x"9C",x"0A",x"CF",x"AB",x"C7",x"DF",x"9C",x"09",x"CF",x"AB",x"C6",x"DF",x"9C",x"08",x"CF",x"A2",x"03",x"BD",x"08",x"CF",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"20",x"77",x"C6",x"20",x"FA",x"C5",x"93",x"90",x"02",x"20",x"AC",x"C6",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"2E",x"2E",x"2E",x"0D",x"00",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"83",x"02",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"7B",x"02",x"AD",x"11",x"DE",x"D3",x"75",x"02",x"A2",x"03",x"BD",x"0E",x"DE",x"9D",x"10",x"CF",x"9D",x"0C",x"CF",x"BD",x"2C",x"DE",x"9D",x"14",x"CF",x"CA",x"10",x"EE",x"A9",x"00",x"8D",x"12",x"CF",x"8D",x"13",x"CF",x"8D",x"0E",x"CF",x"8D",x"0F",x"CF",x"AC",x"10",x"DE",x"F0",x"18",x"A2",x"00",x"18",x"08",x"28",x"BD",x"10",x"CF",x"7D",x"24",x"DE",x"9D",x"10",x"CF",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"88",x"D0",x"E8",x"38",x"A2",x"03",x"BD",x"20",x"DE",x"FD",x"10",x"CF",x"9D",x"1C",x"CF",x"9D",x"20",x"CF",x"CA",x"10",x"F1",x"AD",x"0D",x"DE",x"8D",x"24",x"CF",x"A8",x"29",x"FE",x"F0",x"14",x"A2",x"03",x"18",x"BD",x"20",x"CF",x"6A",x"9D",x"20",x"CF",x"CA",x"10",x"F6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"AD",x"23",x"CF",x"0D",x"22",x"CF",x"F3",x"FC",x"01",x"A2",x"03",x"BD",x"2C",x"DE",x"9D",x"18",x"CF",x"9D",x"4A",x"CF",x"CA",x"10",x"F4",x"20",x"AC",x"C6",x"53",x"45",x"41",x"52",x"43",x"48",x"49",x"4E",x"47",x"20",x"44",x"49",x"52",x"45",x"43",x"54",x"4F",x"52",x"59",x"2E",x"2E",x"2E",x"0D",x"00",x"A9",x"00",x"8D",x"8B",x"D6",x"20",x"78",x"C3",x"20",x"87",x"C3",x"93",x"B0",x"01",x"EA",x"20",x"9C",x"C3",x"93",x"79",x"01",x"A2",x"00",x"AD",x"31",x"CF",x"20",x"6D",x"C3",x"C9",x"44",x"D0",x"ED",x"AD",x"32",x"CF",x"20",x"6D",x"C3",x"C9",x"38",x"D0",x"E3",x"AD",x"33",x"CF",x"20",x"6D",x"C3",x"C9",x"31",x"D0",x"D9",x"20",x"AC",x"C6",x"4D",x"4F",x"55",x"4E",x"54",x"20",x"00",x"20",x"F3",x"C5",x"A2",x"00",x"BD",x"29",x"CF",x"DA",x"20",x"D2",x"FF",x"FA",x"E8",x"E0",x"08",x"D0",x"F3",x"20",x"AC",x"C6",x"3F",x"20",x"00",x"20",x"F3",x"C5",x"58",x"20",x"E4",x"FF",x"C9",x"00",x"F0",x"F9",x"48",x"A9",x"0D",x"20",x"D2",x"FF",x"78",x"20",x"EC",x"C5",x"68",x"C9",x"59",x"D0",x"9D",x"20",x"EB",x"C3",x"20",x"EE",x"C4",x"20",x"77",x"C6",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"8C",x"D6",x"CA",x"10",x"F7",x"20",x"EB",x"C3",x"A2",x"03",x"BD",x"4A",x"CF",x"9D",x"4F",x"CF",x"CA",x"10",x"F7",x"A9",x"00",x"8D",x"55",x"CF",x"8D",x"56",x"CF",x"A9",x"40",x"8D",x"53",x"CF",x"A9",x"06",x"8D",x"54",x"CF",x"AB",x"24",x"CF",x"6B",x"29",x"01",x"D0",x"0C",x"6B",x"4A",x"4B",x"4E",x"54",x"CF",x"6E",x"53",x"CF",x"4C",x"06",x"C2",x"A2",x"03",x"BD",x"4F",x"CF",x"DD",x"4A",x"CF",x"D3",x"81",x"00",x"CA",x"10",x"F4",x"EE",x"55",x"CF",x"D0",x"03",x"EE",x"56",x"CF",x"18",x"AD",x"4F",x"CF",x"69",x"01",x"8D",x"4F",x"CF",x"AD",x"50",x"CF",x"69",x"00",x"8D",x"50",x"CF",x"AD",x"51",x"CF",x"69",x"00",x"8D",x"51",x"CF",x"AD",x"52",x"CF",x"69",x"00",x"8D",x"52",x"CF",x"20",x"38",x"C4",x"B0",x"C4",x"AD",x"53",x"CF",x"CD",x"55",x"CF",x"D0",x"25",x"AD",x"54",x"CF",x"CD",x"56",x"CF",x"D0",x"1D",x"A9",x"07",x"8D",x"8B",x"D6",x"18",x"20",x"DC",x"C6",x"20",x"AC",x"C6",x"44",x"49",x"53",x"4B",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"2E",x"44",x"38",x"31",x"20",x"46",x"49",x"4C",x"45",x"20",x"48",x"41",x"53",x"20",x"57",x"52",x"4F",x"4E",x"47",x"20",x"4C",x"45",x"4E",x"47",x"54",x"48",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"54",x"48",x"41",x"54",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"20",x"49",x"53",x"20",x"46",x"52",x"41",x"47",x"4D",x"45",x"4E",x"54",x"45",x"44",x"2E",x"0D",x"44",x"45",x"2D",x"46",x"52",x"41",x"47",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"20",x"42",x"45",x"46",x"4F",x"52",x"45",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"4E",x"4F",x"20",x"4D",x"4F",x"52",x"45",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"53",x"2E",x"20",x"44",x"52",x"49",x"56",x"45",x"20",x"4D",x"41",x"52",x"4B",x"45",x"44",x"20",x"45",x"4D",x"50",x"54",x"59",x"2E",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"53",x"44",x"2D",x"43",x"41",x"52",x"44",x"20",x"45",x"52",x"52",x"4F",x"52",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"49",x"4E",x"56",x"41",x"4C",x"49",x"44",x"20",x"4F",x"52",x"20",x"55",x"4E",x"53",x"55",x"50",x"50",x"4F",x"52",x"54",x"45",x"44",x"20",x"46",x"49",x"4C",x"45",x"20",x"53",x"59",x"53",x"54",x"45",x"4D",x"2E",x"0D",x"28",x"53",x"48",x"4F",x"55",x"4C",x"44",x"20",x"42",x"45",x"20",x"46",x"41",x"54",x"33",x"32",x"29",x"0D",x"00",x"4C",x"EF",x"C6",x"C9",x"60",x"90",x"06",x"C9",x"7A",x"B0",x"02",x"29",x"5F",x"60",x"A2",x"00",x"BD",x"18",x"CF",x"9D",x"25",x"CF",x"E8",x"E0",x"04",x"D0",x"F5",x"38",x"60",x"A2",x"00",x"BD",x"25",x"CF",x"9D",x"4A",x"CF",x"E8",x"E0",x"04",x"D0",x"F5",x"A9",x"00",x"8D",x"49",x"CF",x"4C",x"05",x"C4",x"AD",x"49",x"CF",x"C9",x"10",x"90",x"0B",x"A9",x"00",x"8D",x"49",x"CF",x"20",x"16",x"C4",x"B0",x"01",x"60",x"A0",x"00",x"AD",x"49",x"CF",x"29",x"08",x"D0",x"1A",x"AD",x"49",x"CF",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DE",x"99",x"29",x"CF",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CF",x"38",x"60",x"AD",x"49",x"CF",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DF",x"99",x"29",x"CF",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CF",x"38",x"60",x"AD",x"3D",x"CF",x"8D",x"4C",x"CF",x"AD",x"3E",x"CF",x"8D",x"4D",x"CF",x"AD",x"43",x"CF",x"8D",x"4A",x"CF",x"AD",x"44",x"CF",x"8D",x"4B",x"CF",x"38",x"60",x"A9",x"00",x"8D",x"4E",x"CF",x"20",x"EE",x"C4",x"B0",x"01",x"60",x"20",x"77",x"C6",x"4C",x"FA",x"C5",x"20",x"43",x"C6",x"EE",x"4E",x"CF",x"AD",x"4E",x"CF",x"CD",x"24",x"CF",x"D0",x"11",x"A9",x"00",x"8D",x"4E",x"CF",x"20",x"38",x"C4",x"B0",x"01",x"60",x"20",x"EE",x"C4",x"20",x"77",x"C6",x"4C",x"FA",x"C5",x"A2",x"00",x"BD",x"4A",x"CF",x"9D",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F5",x"A0",x"07",x"18",x"6E",x"84",x"D6",x"6E",x"83",x"D6",x"6E",x"82",x"D6",x"6E",x"81",x"D6",x"88",x"D0",x"F0",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"0C",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"20",x"77",x"C6",x"20",x"FA",x"C5",x"90",x"63",x"AD",x"4A",x"CF",x"0A",x"0A",x"AA",x"A0",x"00",x"AD",x"4A",x"CF",x"29",x"40",x"D0",x"0E",x"BD",x"00",x"DE",x"99",x"4A",x"CF",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"80",x"0C",x"BD",x"00",x"DF",x"99",x"4A",x"CF",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"AD",x"4D",x"CF",x"29",x"0F",x"8D",x"4D",x"CF",x"AD",x"4D",x"CF",x"0D",x"4C",x"CF",x"0D",x"4B",x"CF",x"0D",x"4A",x"CF",x"C9",x"00",x"F0",x"22",x"AD",x"4D",x"CF",x"C9",x"0F",x"D0",x"19",x"AD",x"4C",x"CF",x"C9",x"FF",x"D0",x"12",x"AD",x"4B",x"CF",x"C9",x"FF",x"D0",x"0B",x"AD",x"4A",x"CF",x"C9",x"FF",x"F0",x"06",x"C9",x"F7",x"F0",x"02",x"38",x"60",x"18",x"60",x"A2",x"03",x"BD",x"4A",x"CF",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A2",x"03",x"38",x"08",x"28",x"BD",x"81",x"D6",x"FD",x"14",x"CF",x"9D",x"81",x"D6",x"08",x"CA",x"10",x"F2",x"28",x"AD",x"24",x"CF",x"A8",x"29",x"FE",x"F0",x"14",x"18",x"2E",x"81",x"D6",x"2E",x"82",x"D6",x"2E",x"83",x"D6",x"2E",x"84",x"D6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"A2",x"00",x"BD",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"10",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CF",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"38",x"60",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"4C",x"FA",x"C5",x"A9",x"42",x"8D",x"80",x"D6",x"A9",x"00",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F9",x"60",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F9",x"60",x"20",x"AF",x"C5",x"20",x"EC",x"C5",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"AD",x"80",x"D6",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F6",x"60",x"38",x"60",x"20",x"C2",x"C5",x"EE",x"57",x"CF",x"D0",x"FB",x"EE",x"58",x"CF",x"D0",x"F6",x"EE",x"59",x"CF",x"D0",x"F1",x"60",x"A9",x"00",x"8D",x"57",x"CF",x"8D",x"58",x"CF",x"A9",x"E0",x"8D",x"59",x"CF",x"60",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"13",x"EE",x"57",x"CF",x"D0",x"0C",x"EE",x"58",x"CF",x"D0",x"07",x"EE",x"59",x"CF",x"D0",x"02",x"A9",x"00",x"18",x"60",x"38",x"60",x"A9",x"81",x"8D",x"80",x"D6",x"38",x"60",x"A9",x"82",x"8D",x"80",x"D6",x"38",x"60",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"40",x"4C",x"16",x"C6",x"EE",x"20",x"D0",x"A2",x"F0",x"A0",x"00",x"A3",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"E8",x"D0",x"F7",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"05",x"D0",x"F9",x"4C",x"3B",x"C6",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"EF",x"AD",x"88",x"D6",x"AD",x"89",x"D6",x"C9",x"02",x"D0",x"CB",x"38",x"60",x"20",x"6F",x"C5",x"4C",x"16",x"C6",x"18",x"60",x"AD",x"80",x"D6",x"29",x"10",x"D0",x"1A",x"AD",x"82",x"D6",x"18",x"69",x"02",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"69",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"69",x"00",x"8D",x"84",x"D6",x"60",x"EE",x"81",x"D6",x"90",x"0D",x"EE",x"82",x"D6",x"90",x"08",x"EE",x"83",x"D6",x"90",x"03",x"EE",x"84",x"D6",x"60",x"AD",x"80",x"D6",x"29",x"10",x"F0",x"01",x"60",x"AD",x"83",x"D6",x"8D",x"84",x"D6",x"AD",x"82",x"D6",x"8D",x"83",x"D6",x"AD",x"81",x"D6",x"8D",x"82",x"D6",x"A9",x"00",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"0A",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"2A",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"2A",x"8D",x"84",x"D6",x"60",x"20",x"F3",x"C5",x"58",x"68",x"8D",x"BB",x"C6",x"68",x"8D",x"BC",x"C6",x"A2",x"01",x"BD",x"FF",x"FF",x"F0",x"06",x"20",x"D2",x"FF",x"E8",x"D0",x"F5",x"38",x"8A",x"6D",x"BB",x"C6",x"8D",x"DA",x"C6",x"A9",x"00",x"6D",x"BC",x"C6",x"8D",x"DB",x"C6",x"78",x"20",x"EC",x"C5",x"4C",x"FF",x"FF",x"B0",x"06",x"A9",x"00",x"8D",x"2F",x"D0",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"60",x"20",x"F3",x"C5",x"18",x"20",x"DC",x"C6",x"AE",x"5A",x"CF",x"9A",x"A9",x"00",x"58",x"18",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"CF",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"A9",x"FF",x"A2",x"0F",x"A0",x"00",x"A3",x"00",x"5C",x"EA",x"A9",x"80",x"A2",x"8D",x"A0",x"00",x"A3",x"00",x"5C",x"EA",x"AD",x"E1",x"D6",x"4A",x"29",x"02",x"09",x"01",x"8D",x"E1",x"D6",x"AD",x"E1",x"D6",x"29",x"20",x"F0",x"F9",x"AD",x"E1",x"D6",x"29",x"04",x"4A",x"09",x"01",x"8D",x"E1",x"D6",x"AD",x"10",x"68",x"C9",x"45",x"D0",x"E7",x"AD",x"19",x"68",x"C9",x"11",x"D0",x"E0",x"AD",x"26",x"68",x"C9",x"11",x"D0",x"D9",x"AD",x"27",x"68",x"C9",x"9E",x"D0",x"D2",x"AD",x"2C",x"68",x"C9",x"A9",x"D0",x"CB",x"20",x"2C",x"68",x"4C",x"A9",x"CF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

begin

--process for read and write operation.
  PROCESS(Clk,cs,ram,address)
  BEGIN
    if(rising_edge(Clk)) then 
      if cs='1' then
        if(we='1') then
          ram(to_integer(unsigned(address))) <= data_i;
        end if;
        data_o <= ram(to_integer(unsigned(address)));
      end if;
    end if;
    if cs='1' then
      data_o <= ram(to_integer(unsigned(address)));
    else
      data_o <= "ZZZZZZZZ";
    end if;
  END PROCESS;

end Behavioral;
