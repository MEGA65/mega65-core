library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

--
entity kickstart is
  port (Clk : in std_logic;
        address : in std_logic_vector(13 downto 0);
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        we : in std_logic;
        -- chip select, active low       
        cs : in std_logic;
        data_i : in std_logic_vector(7 downto 0);
        data_o : out std_logic_vector(7 downto 0)
        );
end kickstart;

architecture Behavioral of kickstart is

-- 16K x 8bit pre-initialised RAM
  type ram_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal ram : ram_t := (x"4C",x"2F",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"39",x"8C",x"EA",x"4C",x"1B",x"8B",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"4C",x"03",x"82",x"EA",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4C",x"42",x"8C",x"AD",x"47",x"D6",x"29",x"FE",x"8D",x"47",x"D6",x"A9",x"FF",x"8D",x"40",x"D6",x"8D",x"7F",x"D6",x"AD",x"47",x"D6",x"09",x"01",x"8D",x"47",x"D6",x"8D",x"7F",x"D6",x"8D",x"40",x"D6",x"AD",x"47",x"D6",x"09",x"01",x"8D",x"47",x"D6",x"8D",x"7F",x"D6",x"4C",x"03",x"82",x"8A",x"29",x"FE",x"30",x"F8",x"AA",x"7C",x"38",x"82",x"A8",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"2C",x"82",x"2C",x"82",x"2C",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"BF",x"82",x"A9",x"01",x"8D",x"41",x"D6",x"A9",x"01",x"8D",x"40",x"D6",x"A9",x"01",x"8D",x"43",x"D6",x"A9",x"01",x"8D",x"42",x"D6",x"4C",x"13",x"82",x"4C",x"2C",x"82",x"A9",x"FF",x"8D",x"80",x"BD",x"8D",x"A0",x"BD",x"8D",x"C0",x"BD",x"8D",x"E0",x"BD",x"38",x"60",x"A9",x"00",x"8D",x"F9",x"BC",x"20",x"49",x"83",x"20",x"35",x"83",x"93",x"BA",x"00",x"20",x"33",x"90",x"A9",x"02",x"8D",x"F9",x"BC",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"AA",x"00",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"A2",x"00",x"A9",x"BE",x"8D",x"01",x"BF",x"A9",x"DF",x"8D",x"02",x"BF",x"20",x"4F",x"83",x"20",x"35",x"83",x"93",x"8F",x"00",x"A9",x"CE",x"8D",x"01",x"BF",x"20",x"4F",x"83",x"20",x"35",x"83",x"93",x"81",x"00",x"A9",x"DE",x"8D",x"01",x"BF",x"20",x"4F",x"83",x"20",x"35",x"83",x"90",x"73",x"A9",x"EE",x"8D",x"01",x"BF",x"20",x"4F",x"83",x"A9",x"00",x"8D",x"F9",x"BC",x"38",x"60",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"20",x"41",x"90",x"90",x"51",x"60",x"A9",x"00",x"8D",x"01",x"BC",x"60",x"A9",x"00",x"8D",x"F9",x"BC",x"A0",x"04",x"B1",x"01",x"C9",x"0C",x"F0",x"0C",x"C9",x"0B",x"F0",x"08",x"A9",x"01",x"8D",x"F9",x"BC",x"4C",x"97",x"83",x"AD",x"01",x"BC",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"A0",x"08",x"B1",x"01",x"9D",x"00",x"BB",x"E8",x"C8",x"C0",x"10",x"D0",x"F5",x"AD",x"01",x"BC",x"20",x"9B",x"83",x"90",x"13",x"AD",x"01",x"BC",x"F0",x"06",x"A0",x"00",x"B1",x"01",x"10",x"06",x"AD",x"01",x"BC",x"8D",x"02",x"BC",x"38",x"60",x"18",x"60",x"A9",x"00",x"8D",x"F9",x"BC",x"0A",x"0A",x"0A",x"0A",x"0A",x"8D",x"04",x"BC",x"09",x"00",x"A8",x"A2",x"00",x"B9",x"00",x"BB",x"9D",x"81",x"D6",x"C8",x"E8",x"E0",x"04",x"D0",x"F4",x"20",x"E2",x"90",x"20",x"41",x"90",x"90",x"D8",x"20",x"33",x"90",x"A9",x"02",x"8D",x"F9",x"BC",x"AD",x"FE",x"DF",x"C9",x"55",x"D0",x"C9",x"AD",x"FF",x"DF",x"C9",x"AA",x"D0",x"C2",x"A9",x"03",x"8D",x"F9",x"BC",x"AD",x"11",x"DE",x"D0",x"B8",x"AD",x"04",x"BC",x"09",x"17",x"A8",x"AD",x"10",x"DE",x"99",x"00",x"BB",x"AD",x"04",x"BC",x"09",x"0D",x"A8",x"A2",x"00",x"BD",x"0E",x"DE",x"99",x"00",x"BB",x"C8",x"E8",x"E0",x"02",x"D0",x"F4",x"AD",x"04",x"BC",x"09",x"09",x"A8",x"A2",x"00",x"BD",x"24",x"DE",x"99",x"00",x"BB",x"C8",x"E8",x"E0",x"04",x"D0",x"F4",x"A9",x"04",x"8D",x"F9",x"BC",x"AD",x"2D",x"DE",x"0D",x"2E",x"DE",x"0D",x"2F",x"DE",x"F0",x"03",x"4C",x"99",x"83",x"AC",x"04",x"BC",x"AD",x"2C",x"DE",x"99",x"0F",x"BB",x"AD",x"04",x"BC",x"09",x"0D",x"A8",x"AD",x"04",x"BC",x"09",x"18",x"AA",x"A3",x"02",x"B9",x"00",x"BB",x"9D",x"00",x"BB",x"C8",x"E8",x"3B",x"D0",x"F5",x"6B",x"9D",x"00",x"BB",x"9D",x"01",x"BB",x"A9",x"05",x"8D",x"F9",x"BC",x"AB",x"10",x"DE",x"F3",x"3E",x"FF",x"C2",x"02",x"D3",x"39",x"FF",x"AD",x"04",x"BC",x"09",x"18",x"A8",x"A2",x"00",x"18",x"08",x"28",x"B9",x"00",x"BB",x"7D",x"24",x"DE",x"99",x"00",x"BB",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"3B",x"D0",x"E1",x"AD",x"04",x"BC",x"09",x"18",x"AA",x"AD",x"04",x"BC",x"09",x"12",x"A8",x"38",x"AD",x"20",x"DE",x"FD",x"00",x"BB",x"99",x"00",x"BB",x"AD",x"21",x"DE",x"FD",x"01",x"BB",x"99",x"01",x"BB",x"AD",x"22",x"DE",x"FD",x"02",x"BB",x"99",x"02",x"BB",x"AD",x"23",x"DE",x"FD",x"03",x"BB",x"99",x"03",x"BB",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"AD",x"0D",x"DE",x"99",x"00",x"BB",x"4B",x"29",x"FE",x"F0",x"1E",x"AD",x"04",x"BC",x"09",x"12",x"18",x"69",x"03",x"A8",x"A2",x"03",x"18",x"B9",x"00",x"BB",x"6A",x"99",x"00",x"BB",x"88",x"CA",x"10",x"F5",x"6B",x"4A",x"4B",x"29",x"FE",x"D0",x"E2",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"AD",x"0D",x"DE",x"99",x"00",x"BB",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"A9",x"06",x"8D",x"F9",x"BC",x"B9",x"03",x"BB",x"19",x"02",x"BB",x"F3",x"9A",x"FE",x"AD",x"04",x"BC",x"09",x"10",x"A8",x"A2",x"03",x"BD",x"2C",x"DE",x"99",x"00",x"BB",x"CA",x"10",x"F7",x"AD",x"04",x"BC",x"09",x"08",x"A8",x"A9",x"0F",x"99",x"00",x"BB",x"EE",x"01",x"BC",x"A9",x"00",x"8D",x"F9",x"BC",x"38",x"60",x"8D",x"F9",x"BC",x"18",x"60",x"A9",x"80",x"EC",x"01",x"BC",x"B3",x"67",x"FE",x"8E",x"03",x"BC",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8D",x"04",x"BC",x"38",x"60",x"20",x"2B",x"85",x"90",x"E3",x"AE",x"04",x"BC",x"BD",x"10",x"BB",x"8D",x"05",x"BC",x"BD",x"11",x"BB",x"8D",x"06",x"BC",x"A9",x"00",x"8D",x"07",x"BC",x"8D",x"08",x"BC",x"4C",x"1F",x"85",x"A2",x"03",x"BD",x"B2",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"AD",x"81",x"D6",x"38",x"E9",x"02",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"E9",x"00",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"E9",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"E9",x"00",x"8D",x"84",x"D6",x"AE",x"04",x"BC",x"BD",x"16",x"BB",x"A8",x"29",x"FE",x"F0",x"14",x"18",x"2E",x"81",x"D6",x"2E",x"82",x"D6",x"2E",x"83",x"D6",x"2E",x"84",x"D6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"A2",x"00",x"BD",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F8",x"AD",x"04",x"BC",x"09",x"18",x"A8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"79",x"00",x"BB",x"9D",x"81",x"D6",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"AD",x"04",x"BC",x"09",x"00",x"A8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"79",x"00",x"BB",x"9D",x"81",x"D6",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"38",x"60",x"AE",x"69",x"BC",x"E0",x"3F",x"A9",x"81",x"B3",x"2E",x"FF",x"BD",x"6A",x"BC",x"20",x"84",x"8F",x"9D",x"6A",x"BC",x"E8",x"EC",x"69",x"BC",x"D0",x"F1",x"38",x"60",x"A2",x"00",x"8A",x"0A",x"0A",x"0A",x"0A",x"A8",x"B9",x"B7",x"BC",x"C9",x"FF",x"F0",x"0A",x"E8",x"E0",x"04",x"D0",x"EE",x"A9",x"84",x"4C",x"26",x"85",x"A0",x"0F",x"A9",x"00",x"99",x"B7",x"BC",x"88",x"D0",x"FA",x"8E",x"F7",x"BC",x"8A",x"0A",x"0A",x"0A",x"0A",x"8D",x"F8",x"BC",x"38",x"60",x"A9",x"FF",x"8D",x"B7",x"BC",x"8D",x"C7",x"BC",x"8D",x"D7",x"BC",x"8D",x"E7",x"BC",x"38",x"60",x"AE",x"F8",x"BC",x"BD",x"B8",x"BC",x"C9",x"01",x"D0",x"00",x"AE",x"F8",x"BC",x"A9",x"FF",x"9D",x"B7",x"BC",x"38",x"60",x"AD",x"68",x"BC",x"29",x"10",x"F0",x"05",x"A9",x"86",x"4C",x"26",x"85",x"20",x"97",x"88",x"93",x"BA",x"FE",x"4C",x"CF",x"88",x"20",x"80",x"86",x"08",x"20",x"4A",x"86",x"28",x"93",x"AC",x"FE",x"38",x"60",x"20",x"EF",x"85",x"93",x"A4",x"FE",x"20",x"A3",x"86",x"93",x"9E",x"FE",x"4C",x"8F",x"86",x"20",x"D5",x"86",x"B0",x"08",x"20",x"4A",x"86",x"A9",x"88",x"4C",x"26",x"85",x"20",x"58",x"88",x"90",x"EE",x"38",x"60",x"20",x"0A",x"86",x"93",x"81",x"FE",x"8A",x"0A",x"0A",x"0A",x"0A",x"A8",x"AD",x"03",x"BC",x"99",x"B7",x"BC",x"A2",x"00",x"BD",x"05",x"BC",x"99",x"B9",x"BC",x"99",x"BD",x"BC",x"C8",x"E8",x"E0",x"04",x"D0",x"F1",x"AE",x"F8",x"BC",x"A9",x"80",x"9D",x"B8",x"BC",x"20",x"CF",x"88",x"93",x"56",x"FE",x"60",x"A9",x"00",x"8D",x"52",x"BC",x"20",x"0C",x"89",x"AE",x"F8",x"BC",x"BD",x"B8",x"BC",x"C9",x"80",x"F0",x"0E",x"C9",x"81",x"D0",x"05",x"A9",x"FF",x"4C",x"26",x"85",x"A9",x"87",x"4C",x"26",x"85",x"A2",x"54",x"A9",x"00",x"9D",x"0F",x"BC",x"CA",x"10",x"FA",x"20",x"0C",x"89",x"93",x"25",x"FE",x"20",x"33",x"90",x"AD",x"F8",x"BC",x"09",x"0B",x"AA",x"BD",x"B7",x"BC",x"8D",x"01",x"BF",x"BD",x"B8",x"BC",x"18",x"69",x"DE",x"8D",x"02",x"BF",x"A0",x"0B",x"B1",x"01",x"C9",x"0F",x"D3",x"72",x"00",x"A0",x"0C",x"B1",x"01",x"D3",x"6B",x"00",x"A9",x"00",x"29",x"3F",x"C9",x"04",x"B0",x"55",x"AA",x"BD",x"53",x"88",x"AA",x"A0",x"01",x"A3",x"05",x"B1",x"01",x"F0",x"37",x"9D",x"0F",x"BC",x"E8",x"E0",x"40",x"F0",x"2F",x"C8",x"C8",x"3B",x"D0",x"EF",x"A0",x"0E",x"A3",x"06",x"B1",x"01",x"F0",x"22",x"9D",x"0F",x"BC",x"E8",x"E0",x"40",x"F0",x"1A",x"C8",x"C8",x"3B",x"D0",x"EF",x"A0",x"1C",x"A3",x"02",x"B1",x"01",x"F0",x"0D",x"9D",x"0F",x"BC",x"E8",x"E0",x"40",x"F0",x"05",x"C8",x"C8",x"3B",x"D0",x"EF",x"EC",x"52",x"BC",x"90",x"0C",x"8E",x"52",x"BC",x"E0",x"3F",x"B0",x"05",x"A9",x"00",x"9D",x"0F",x"BC",x"20",x"73",x"88",x"90",x"03",x"4C",x"08",x"87",x"A9",x"FF",x"4C",x"26",x"85",x"A0",x"00",x"B1",x"01",x"F3",x"AD",x"00",x"C9",x"E5",x"F3",x"A8",x"00",x"A2",x"00",x"B1",x"01",x"9D",x"53",x"BC",x"E8",x"C8",x"E0",x"0B",x"D0",x"F5",x"AD",x"52",x"BC",x"D0",x"3B",x"A0",x"00",x"A2",x"00",x"B1",x"01",x"9D",x"0F",x"BC",x"E8",x"C8",x"C9",x"20",x"F0",x"05",x"E0",x"08",x"D0",x"F1",x"E8",x"CA",x"A9",x"2E",x"9D",x"0F",x"BC",x"E8",x"A0",x"08",x"A3",x"00",x"B1",x"01",x"9D",x"0F",x"BC",x"E8",x"C8",x"1B",x"C2",x"03",x"F0",x"08",x"C9",x"20",x"F0",x"04",x"E0",x"0C",x"D0",x"EC",x"A9",x"00",x"9D",x"0F",x"BC",x"8E",x"52",x"BC",x"A0",x"1A",x"B1",x"01",x"8D",x"60",x"BC",x"C8",x"B1",x"01",x"8D",x"61",x"BC",x"A0",x"14",x"B1",x"01",x"8D",x"62",x"BC",x"C8",x"B1",x"01",x"8D",x"63",x"BC",x"A0",x"1C",x"A2",x"00",x"B1",x"01",x"9D",x"64",x"BC",x"C8",x"E8",x"E0",x"04",x"D0",x"F5",x"A0",x"0B",x"B1",x"01",x"8D",x"68",x"BC",x"20",x"73",x"88",x"B0",x"0E",x"AE",x"F8",x"BC",x"A9",x"81",x"9D",x"B8",x"BC",x"AE",x"F8",x"BC",x"BD",x"B8",x"BC",x"AD",x"52",x"BC",x"C9",x"00",x"F3",x"9B",x"FE",x"AD",x"53",x"BC",x"C9",x"20",x"F3",x"93",x"FE",x"C9",x"00",x"F3",x"8E",x"FE",x"38",x"60",x"20",x"73",x"88",x"B3",x"86",x"FE",x"4C",x"29",x"85",x"00",x"0E",x"1C",x"2A",x"38",x"AD",x"52",x"BC",x"CD",x"69",x"BC",x"D0",x"11",x"AE",x"52",x"BC",x"CA",x"BD",x"0F",x"BC",x"DD",x"6A",x"BC",x"D0",x"05",x"CA",x"D0",x"F5",x"38",x"60",x"18",x"60",x"AC",x"F8",x"BC",x"18",x"B9",x"C2",x"BC",x"69",x"20",x"99",x"C2",x"BC",x"D0",x"0B",x"B9",x"C3",x"BC",x"1A",x"C9",x"01",x"D0",x"05",x"99",x"C3",x"BC",x"38",x"60",x"A9",x"00",x"99",x"C3",x"BC",x"20",x"35",x"89",x"60",x"20",x"0A",x"86",x"20",x"F1",x"88",x"AD",x"03",x"BC",x"9D",x"B7",x"BC",x"A0",x"00",x"B9",x"60",x"BC",x"9D",x"B9",x"BC",x"9D",x"BD",x"BC",x"E8",x"C8",x"C0",x"04",x"D0",x"F1",x"20",x"F1",x"88",x"AD",x"03",x"BC",x"9D",x"B7",x"BC",x"A9",x"00",x"9D",x"B8",x"BC",x"A9",x"00",x"9D",x"C1",x"BC",x"9D",x"C2",x"BC",x"9D",x"C3",x"BC",x"38",x"60",x"20",x"F1",x"88",x"A0",x"03",x"BD",x"B9",x"BC",x"9D",x"BD",x"BC",x"E8",x"88",x"10",x"F6",x"20",x"F1",x"88",x"A9",x"00",x"A0",x"06",x"9D",x"C1",x"BC",x"E8",x"88",x"D0",x"F9",x"20",x"F1",x"88",x"38",x"60",x"AD",x"F7",x"BC",x"0A",x"0A",x"0A",x"0A",x"AA",x"60",x"20",x"F1",x"88",x"A0",x"00",x"BD",x"BD",x"BC",x"99",x"B2",x"BC",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"60",x"20",x"FA",x"88",x"20",x"60",x"85",x"20",x"F1",x"88",x"09",x"0A",x"A8",x"A2",x"00",x"18",x"B9",x"B7",x"BC",x"D0",x"02",x"A9",x"00",x"7D",x"81",x"D6",x"9D",x"81",x"D6",x"90",x"05",x"E8",x"E0",x"04",x"D0",x"F1",x"20",x"E2",x"90",x"4C",x"41",x"90",x"AE",x"F8",x"BC",x"BD",x"C4",x"BC",x"18",x"69",x"02",x"9D",x"C4",x"BC",x"90",x"08",x"FE",x"C5",x"BC",x"D0",x"03",x"FE",x"C6",x"BC",x"FE",x"C1",x"BC",x"BD",x"C1",x"BC",x"AC",x"04",x"BC",x"D9",x"16",x"BB",x"F0",x"02",x"38",x"60",x"AC",x"F8",x"BC",x"A9",x"00",x"99",x"C1",x"BC",x"20",x"FA",x"88",x"A2",x"03",x"BD",x"B2",x"BC",x"9D",x"AE",x"BC",x"CA",x"10",x"F7",x"AD",x"B2",x"BC",x"8D",x"05",x"BF",x"A0",x"07",x"18",x"6E",x"B5",x"BC",x"6E",x"B4",x"BC",x"6E",x"B3",x"BC",x"6E",x"B2",x"BC",x"88",x"D0",x"F0",x"AC",x"04",x"BC",x"A2",x"00",x"18",x"08",x"28",x"BD",x"B2",x"BC",x"79",x"00",x"BB",x"9D",x"B2",x"BC",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"AC",x"04",x"BC",x"A2",x"00",x"18",x"08",x"28",x"BD",x"B2",x"BC",x"79",x"0D",x"BB",x"9D",x"B2",x"BC",x"08",x"C8",x"E8",x"E0",x"02",x"D0",x"EF",x"A2",x"03",x"BD",x"B2",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"28",x"BD",x"B2",x"BC",x"69",x"00",x"9D",x"B2",x"BC",x"08",x"E8",x"E0",x"04",x"D0",x"F1",x"28",x"20",x"E2",x"90",x"20",x"41",x"90",x"93",x"4C",x"FB",x"20",x"33",x"90",x"AD",x"05",x"BF",x"0A",x"0A",x"AA",x"AD",x"F8",x"BC",x"09",x"06",x"A8",x"8C",x"06",x"BF",x"AC",x"06",x"BF",x"A3",x"00",x"AD",x"05",x"BF",x"29",x"40",x"D0",x"0F",x"BD",x"00",x"DE",x"99",x"B7",x"BC",x"E8",x"C8",x"1B",x"C2",x"04",x"D0",x"F3",x"80",x"0D",x"BD",x"00",x"DF",x"99",x"B7",x"BC",x"E8",x"C8",x"1B",x"C2",x"04",x"D0",x"F3",x"A0",x"00",x"B9",x"BA",x"BC",x"4B",x"5A",x"20",x"AD",x"94",x"7A",x"B9",x"B9",x"BC",x"4B",x"5A",x"20",x"AD",x"94",x"7A",x"B9",x"B8",x"BC",x"4B",x"5A",x"20",x"AD",x"94",x"7A",x"B9",x"B7",x"BC",x"4B",x"20",x"AD",x"94",x"AC",x"06",x"BF",x"B9",x"BA",x"BC",x"29",x"0F",x"99",x"BA",x"BC",x"B9",x"BA",x"BC",x"19",x"B9",x"BC",x"19",x"B8",x"BC",x"19",x"B7",x"BC",x"C9",x"00",x"F0",x"22",x"B9",x"BA",x"BC",x"C9",x"0F",x"D0",x"19",x"B9",x"B9",x"BC",x"C9",x"FF",x"D0",x"12",x"B9",x"B8",x"BC",x"C9",x"FF",x"D0",x"0B",x"B9",x"B7",x"BC",x"C9",x"FF",x"F0",x"06",x"C9",x"F7",x"F0",x"02",x"38",x"60",x"A9",x"85",x"4C",x"26",x"85",x"A2",x"6B",x"A0",x"99",x"20",x"29",x"94",x"A0",x"00",x"AB",x"B5",x"BC",x"20",x"AD",x"94",x"AB",x"B4",x"BC",x"20",x"AD",x"94",x"AB",x"B3",x"BC",x"20",x"AD",x"94",x"AB",x"B2",x"BC",x"4C",x"AD",x"94",x"A2",x"00",x"8E",x"AC",x"BC",x"8E",x"AD",x"BC",x"20",x"80",x"86",x"08",x"20",x"4A",x"86",x"28",x"93",x"78",x"FA",x"20",x"5E",x"86",x"93",x"72",x"FA",x"20",x"33",x"90",x"20",x"0C",x"89",x"90",x"33",x"A2",x"00",x"A3",x"00",x"BD",x"00",x"DE",x"EA",x"92",x"17",x"1B",x"E8",x"D0",x"F6",x"E3",x"18",x"BD",x"00",x"DF",x"EA",x"92",x"17",x"1B",x"E8",x"D0",x"F6",x"20",x"35",x"89",x"90",x"14",x"E3",x"18",x"EE",x"AC",x"BC",x"D0",x"D5",x"EE",x"AD",x"BC",x"D0",x"D0",x"20",x"4A",x"86",x"A9",x"83",x"4C",x"26",x"85",x"20",x"4A",x"86",x"4C",x"1F",x"85",x"8E",x"01",x"BF",x"8C",x"02",x"BF",x"A0",x"00",x"B1",x"01",x"99",x"6A",x"BC",x"F0",x"0E",x"C8",x"C0",x"40",x"D0",x"F4",x"A9",x"00",x"8D",x"69",x"BC",x"A9",x"81",x"18",x"60",x"8C",x"69",x"BC",x"38",x"60",x"20",x"09",x"8C",x"A2",x"4B",x"A0",x"8B",x"20",x"29",x"94",x"A0",x"00",x"AB",x"49",x"D6",x"20",x"AD",x"94",x"AB",x"48",x"D6",x"20",x"AD",x"94",x"AB",x"4F",x"D6",x"20",x"AD",x"94",x"AB",x"4A",x"D6",x"20",x"AD",x"94",x"AB",x"49",x"D6",x"20",x"AD",x"94",x"EE",x"20",x"D0",x"4C",x"45",x"8B",x"50",x"41",x"47",x"45",x"20",x"46",x"41",x"55",x"4C",x"54",x"3A",x"20",x"50",x"43",x"3D",x"24",x"24",x"24",x"24",x"2C",x"20",x"4D",x"41",x"50",x"3D",x"24",x"24",x"2E",x"24",x"24",x"24",x"24",x"2E",x"30",x"30",x"20",x"20",x"20",x"20",x"20",x"A9",x"00",x"60",x"A9",x"00",x"8D",x"40",x"D6",x"8D",x"41",x"D6",x"8D",x"42",x"D6",x"8D",x"43",x"D6",x"8D",x"44",x"D6",x"A9",x"FF",x"8D",x"45",x"D6",x"A9",x"01",x"8D",x"46",x"D6",x"A9",x"F7",x"8D",x"47",x"D6",x"A9",x"00",x"8D",x"4A",x"D6",x"8D",x"4B",x"D6",x"8D",x"4C",x"D6",x"8D",x"4D",x"D6",x"8D",x"4E",x"D6",x"8D",x"4F",x"D6",x"A9",x"3F",x"8D",x"50",x"D6",x"8D",x"51",x"D6",x"A9",x"00",x"8D",x"52",x"D6",x"60",x"A2",x"FC",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"0B",x"95",x"AD",x"00",x"BC",x"8D",x"48",x"D6",x"A2",x"FC",x"E8",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"0B",x"95",x"AD",x"00",x"BC",x"8D",x"49",x"D6",x"60",x"A9",x"00",x"A2",x"5D",x"9D",x"00",x"D6",x"E8",x"E0",x"70",x"D0",x"F8",x"60",x"A2",x"00",x"8A",x"9D",x"00",x"BD",x"E8",x"D0",x"FA",x"20",x"DC",x"8B",x"4C",x"C2",x"82",x"20",x"E9",x"8B",x"20",x"73",x"8B",x"8D",x"00",x"BD",x"60",x"20",x"F8",x"8B",x"20",x"76",x"8B",x"60",x"78",x"D8",x"03",x"A9",x"00",x"8D",x"17",x"D0",x"A9",x"7F",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"A9",x"00",x"8D",x"1A",x"D0",x"A9",x"7F",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"A9",x"00",x"8D",x"19",x"D0",x"38",x"20",x"4D",x"95",x"20",x"D9",x"91",x"20",x"17",x"93",x"20",x"13",x"92",x"60",x"78",x"A9",x"00",x"8D",x"00",x"BF",x"4C",x"4B",x"8C",x"78",x"A9",x"80",x"8D",x"00",x"BF",x"4C",x"4B",x"8C",x"20",x"09",x"8C",x"A2",x"7D",x"A0",x"97",x"20",x"98",x"94",x"A2",x"CA",x"A0",x"9B",x"20",x"29",x"94",x"A2",x"A7",x"A0",x"A7",x"20",x"29",x"94",x"20",x"60",x"95",x"AD",x"00",x"BF",x"30",x"17",x"AD",x"F1",x"D6",x"29",x"02",x"F0",x"10",x"A2",x"1B",x"A0",x"9B",x"20",x"29",x"94",x"20",x"DA",x"95",x"20",x"0C",x"96",x"4C",x"7C",x"8C",x"A2",x"09",x"A0",x"98",x"20",x"29",x"94",x"20",x"8F",x"8F",x"B0",x"03",x"4C",x"89",x"8C",x"20",x"3A",x"86",x"20",x"D2",x"82",x"A2",x"B7",x"A0",x"98",x"20",x"29",x"94",x"A0",x"00",x"AB",x"01",x"BC",x"20",x"AD",x"94",x"AE",x"02",x"BC",x"20",x"41",x"85",x"B0",x"0F",x"A2",x"87",x"A0",x"9B",x"20",x"29",x"94",x"A0",x"00",x"AB",x"F9",x"BC",x"20",x"AD",x"94",x"A9",x"00",x"85",x"17",x"A9",x"40",x"85",x"18",x"A9",x"00",x"85",x"19",x"A9",x"00",x"85",x"1A",x"A2",x"F7",x"A0",x"9B",x"20",x"F9",x"8A",x"20",x"9F",x"8A",x"B0",x"0F",x"A2",x"60",x"A0",x"9B",x"20",x"29",x"94",x"A0",x"00",x"AB",x"F9",x"BC",x"20",x"AD",x"94",x"AD",x"7E",x"D6",x"F0",x"0A",x"A2",x"01",x"A0",x"9B",x"20",x"29",x"94",x"4C",x"7C",x"8D",x"A9",x"00",x"85",x"17",x"A9",x"40",x"85",x"18",x"A9",x"00",x"85",x"19",x"A9",x"00",x"85",x"1A",x"A2",x"EC",x"A0",x"9B",x"20",x"F9",x"8A",x"20",x"9F",x"8A",x"93",x"62",x"00",x"A2",x"DC",x"A0",x"9A",x"20",x"29",x"94",x"A0",x"00",x"AB",x"12",x"00",x"20",x"AD",x"94",x"AB",x"11",x"00",x"20",x"AD",x"94",x"AB",x"10",x"00",x"20",x"AD",x"94",x"AB",x"0F",x"00",x"20",x"AD",x"94",x"A2",x"00",x"BD",x"43",x"8D",x"9D",x"00",x"30",x"E8",x"D0",x"F7",x"4C",x"00",x"30",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"8D",x"06",x"D7",x"A9",x"00",x"8D",x"05",x"D7",x"A9",x"8D",x"8D",x"01",x"D7",x"A9",x"6A",x"8D",x"00",x"D7",x"A9",x"00",x"8D",x"06",x"D7",x"8D",x"7E",x"D6",x"4C",x"00",x"81",x"00",x"00",x"40",x"00",x"40",x"00",x"00",x"80",x"0F",x"00",x"00",x"A2",x"BA",x"A0",x"9A",x"20",x"29",x"94",x"A9",x"00",x"8D",x"8B",x"D6",x"20",x"41",x"85",x"93",x"E4",x"01",x"A2",x"E2",x"A0",x"9B",x"20",x"F9",x"8A",x"20",x"73",x"86",x"93",x"CA",x"00",x"20",x"4A",x"86",x"A2",x"BC",x"A0",x"99",x"20",x"29",x"94",x"20",x"97",x"88",x"93",x"BA",x"00",x"20",x"5E",x"86",x"93",x"B4",x"00",x"A9",x"00",x"8D",x"0E",x"CE",x"8D",x"0F",x"CE",x"A9",x"40",x"8D",x"0C",x"CE",x"A9",x"06",x"8D",x"0D",x"CE",x"AE",x"04",x"BC",x"BD",x"16",x"BB",x"4B",x"6B",x"29",x"01",x"D0",x"0C",x"6B",x"4A",x"4B",x"4E",x"0D",x"CE",x"6E",x"0C",x"CE",x"4C",x"C3",x"8D",x"AE",x"F8",x"BC",x"A0",x"00",x"BD",x"BD",x"BC",x"99",x"08",x"CE",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"AE",x"F8",x"BC",x"A0",x"00",x"BD",x"BD",x"BC",x"D9",x"08",x"CE",x"D3",x"61",x"00",x"E8",x"C8",x"C0",x"04",x"D0",x"F1",x"EE",x"0E",x"CE",x"D0",x"03",x"EE",x"0F",x"CE",x"18",x"AD",x"08",x"CE",x"69",x"01",x"8D",x"08",x"CE",x"AD",x"09",x"CE",x"69",x"00",x"8D",x"09",x"CE",x"AD",x"0A",x"CE",x"69",x"00",x"8D",x"0A",x"CE",x"AD",x"0B",x"CE",x"69",x"00",x"8D",x"0B",x"CE",x"20",x"5B",x"89",x"B0",x"BE",x"20",x"4A",x"86",x"AD",x"0C",x"CE",x"CD",x"0E",x"CE",x"D0",x"17",x"AD",x"0D",x"CE",x"CD",x"0F",x"CE",x"D0",x"0F",x"A9",x"07",x"8D",x"8B",x"D6",x"A2",x"37",x"A0",x"9A",x"20",x"29",x"94",x"4C",x"6C",x"8E",x"A2",x"E5",x"A0",x"99",x"20",x"29",x"94",x"4C",x"6C",x"8E",x"A2",x"0E",x"A0",x"9A",x"20",x"29",x"94",x"4C",x"6C",x"8E",x"A2",x"98",x"A0",x"99",x"20",x"29",x"94",x"A0",x"00",x"AB",x"F9",x"BC",x"20",x"AD",x"94",x"20",x"17",x"91",x"90",x"0A",x"A2",x"94",x"A0",x"97",x"20",x"29",x"94",x"4C",x"D4",x"94",x"A2",x"AE",x"A0",x"97",x"20",x"29",x"94",x"A2",x"CB",x"A0",x"9B",x"20",x"F9",x"8A",x"A9",x"00",x"85",x"17",x"A9",x"E0",x"85",x"18",x"A9",x"F7",x"85",x"19",x"A9",x"0F",x"85",x"1A",x"20",x"9F",x"8A",x"B0",x"0A",x"A2",x"CE",x"A0",x"97",x"20",x"29",x"94",x"4C",x"CC",x"8E",x"AE",x"F8",x"BC",x"BD",x"C4",x"BC",x"8D",x"06",x"CE",x"BD",x"C5",x"BC",x"8D",x"07",x"CE",x"A2",x"E9",x"A0",x"97",x"20",x"29",x"94",x"A0",x"00",x"AB",x"07",x"CE",x"20",x"AD",x"94",x"AB",x"06",x"CE",x"20",x"AD",x"94",x"A2",x"D7",x"A0",x"9B",x"20",x"F9",x"8A",x"A9",x"00",x"85",x"17",x"85",x"18",x"85",x"1A",x"A9",x"02",x"85",x"19",x"20",x"9F",x"8A",x"B0",x"21",x"A2",x"0B",x"BD",x"D7",x"9B",x"9D",x"8B",x"9A",x"CA",x"D0",x"F7",x"A2",x"78",x"A0",x"9A",x"20",x"29",x"94",x"20",x"ED",x"8F",x"20",x"ED",x"8F",x"20",x"ED",x"8F",x"20",x"ED",x"8F",x"4C",x"6A",x"8F",x"AE",x"F8",x"BC",x"BD",x"C4",x"BC",x"8D",x"06",x"CE",x"BD",x"C5",x"BC",x"8D",x"07",x"CE",x"AD",x"06",x"CE",x"D0",x"31",x"AD",x"07",x"CE",x"C9",x"00",x"F0",x"2A",x"C9",x"02",x"D0",x"0D",x"20",x"4A",x"91",x"A2",x"94",x"A0",x"97",x"20",x"29",x"94",x"4C",x"D4",x"94",x"A2",x"2A",x"A0",x"99",x"20",x"29",x"94",x"AB",x"07",x"CE",x"20",x"AD",x"94",x"AB",x"06",x"CE",x"20",x"AD",x"94",x"20",x"ED",x"8F",x"4C",x"39",x"8C",x"A2",x"4A",x"A0",x"99",x"20",x"29",x"94",x"AB",x"07",x"CE",x"20",x"AD",x"94",x"AB",x"06",x"CE",x"20",x"AD",x"94",x"20",x"ED",x"8F",x"4C",x"39",x"8C",x"A2",x"F2",x"A0",x"98",x"20",x"29",x"94",x"A2",x"36",x"A0",x"98",x"20",x"29",x"94",x"20",x"ED",x"8F",x"4C",x"39",x"8C",x"A2",x"51",x"A0",x"98",x"20",x"29",x"94",x"20",x"ED",x"8F",x"4C",x"39",x"8C",x"C9",x"60",x"90",x"06",x"C9",x"7A",x"B0",x"02",x"29",x"5F",x"60",x"20",x"AD",x"8F",x"B0",x"01",x"60",x"A2",x"1F",x"A0",x"98",x"20",x"29",x"94",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"4C",x"41",x"90",x"A9",x"42",x"8D",x"80",x"D6",x"A9",x"00",x"8D",x"80",x"D6",x"20",x"09",x"90",x"20",x"17",x"90",x"B0",x"03",x"D0",x"F9",x"60",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"09",x"90",x"20",x"17",x"90",x"B0",x"03",x"D0",x"F9",x"60",x"20",x"ED",x"8F",x"20",x"33",x"90",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"09",x"90",x"AD",x"80",x"D6",x"20",x"17",x"90",x"B0",x"03",x"D0",x"F6",x"60",x"38",x"60",x"20",x"09",x"90",x"EE",x"20",x"D0",x"20",x"0C",x"96",x"CE",x"20",x"D0",x"EE",x"00",x"03",x"D0",x"F2",x"EE",x"01",x"03",x"D0",x"ED",x"EE",x"02",x"03",x"D0",x"E8",x"60",x"A9",x"00",x"8D",x"00",x"03",x"8D",x"01",x"03",x"A9",x"F7",x"8D",x"02",x"03",x"60",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"13",x"EE",x"00",x"03",x"D0",x"0C",x"EE",x"01",x"03",x"D0",x"07",x"EE",x"02",x"03",x"D0",x"02",x"A9",x"00",x"18",x"60",x"38",x"60",x"A9",x"81",x"8D",x"80",x"D6",x"38",x"60",x"A9",x"82",x"8D",x"80",x"D6",x"38",x"60",x"AD",x"80",x"D6",x"29",x"01",x"D3",x"3E",x"00",x"4C",x"5B",x"90",x"A2",x"F0",x"A0",x"00",x"A3",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"E8",x"D0",x"F7",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"09",x"90",x"20",x"17",x"90",x"B0",x"05",x"D0",x"F9",x"4C",x"80",x"90",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"EF",x"AD",x"88",x"D6",x"AD",x"89",x"D6",x"C9",x"02",x"D0",x"CE",x"38",x"60",x"20",x"AD",x"8F",x"4C",x"5B",x"90",x"A9",x"07",x"8D",x"F9",x"BC",x"18",x"60",x"A2",x"82",x"A0",x"99",x"20",x"29",x"94",x"A0",x"00",x"AB",x"84",x"D6",x"20",x"AD",x"94",x"AB",x"83",x"D6",x"20",x"AD",x"94",x"AB",x"82",x"D6",x"20",x"AD",x"94",x"AB",x"81",x"D6",x"4C",x"AD",x"94",x"AD",x"80",x"D6",x"29",x"10",x"D0",x"1A",x"AD",x"82",x"D6",x"18",x"69",x"02",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"69",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"69",x"00",x"8D",x"84",x"D6",x"60",x"EE",x"81",x"D6",x"90",x"0D",x"EE",x"82",x"D6",x"90",x"08",x"EE",x"83",x"D6",x"90",x"03",x"EE",x"84",x"D6",x"60",x"AD",x"80",x"D6",x"29",x"10",x"F0",x"01",x"60",x"AD",x"83",x"D6",x"8D",x"84",x"D6",x"AD",x"82",x"D6",x"8D",x"83",x"D6",x"AD",x"81",x"D6",x"8D",x"82",x"D6",x"A9",x"00",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"0A",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"2A",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"2A",x"8D",x"84",x"D6",x"60",x"AD",x"F1",x"D6",x"29",x"20",x"D0",x"2A",x"AD",x"DC",x"9B",x"C9",x"2E",x"D0",x"23",x"20",x"74",x"91",x"20",x"60",x"91",x"AD",x"00",x"40",x"CD",x"02",x"CE",x"D0",x"15",x"AD",x"01",x"40",x"CD",x"03",x"CE",x"D0",x"0D",x"AD",x"02",x"40",x"CD",x"04",x"CE",x"D0",x"05",x"20",x"3C",x"95",x"38",x"60",x"18",x"60",x"20",x"60",x"91",x"AD",x"02",x"CE",x"8D",x"00",x"40",x"AD",x"03",x"CE",x"8D",x"01",x"40",x"AD",x"04",x"CE",x"8D",x"02",x"40",x"60",x"A9",x"80",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"A9",x"C0",x"A2",x"CF",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"60",x"A9",x"03",x"8D",x"02",x"CE",x"8D",x"03",x"CE",x"8D",x"04",x"CE",x"8D",x"05",x"CE",x"A9",x"08",x"8D",x"00",x"CE",x"AD",x"00",x"CE",x"38",x"E9",x"01",x"4A",x"4A",x"09",x"C0",x"AA",x"AD",x"00",x"CE",x"38",x"E9",x"01",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A9",x"00",x"85",x"07",x"A9",x"40",x"85",x"08",x"A0",x"00",x"AD",x"02",x"CE",x"18",x"71",x"07",x"8D",x"02",x"CE",x"90",x"08",x"EE",x"03",x"CE",x"90",x"03",x"EE",x"04",x"CE",x"C8",x"D0",x"EA",x"E6",x"08",x"A5",x"08",x"C9",x"80",x"D0",x"E0",x"EE",x"00",x"CE",x"AD",x"00",x"CE",x"C9",x"10",x"D0",x"B1",x"4C",x"3C",x"95",x"A9",x"40",x"8D",x"30",x"D0",x"A9",x"00",x"8D",x"31",x"D0",x"8D",x"20",x"D0",x"8D",x"21",x"D0",x"8D",x"54",x"D0",x"A9",x"14",x"8D",x"18",x"D0",x"A9",x"1B",x"8D",x"11",x"D0",x"A9",x"C8",x"8D",x"16",x"D0",x"A9",x"FF",x"8D",x"01",x"DD",x"8D",x"00",x"DD",x"A9",x"05",x"8D",x"54",x"D0",x"A9",x"50",x"8D",x"40",x"D0",x"A9",x"00",x"8D",x"41",x"D0",x"60",x"A9",x"04",x"8D",x"30",x"D0",x"A9",x"FF",x"8D",x"70",x"D0",x"A9",x"00",x"8D",x"00",x"D1",x"8D",x"00",x"D2",x"8D",x"00",x"D3",x"A9",x"FF",x"8D",x"01",x"D1",x"8D",x"01",x"D2",x"8D",x"01",x"D3",x"A9",x"BA",x"8D",x"02",x"D1",x"A9",x"13",x"8D",x"02",x"D2",x"A9",x"62",x"8D",x"02",x"D3",x"A9",x"66",x"8D",x"03",x"D1",x"A9",x"AD",x"8D",x"03",x"D2",x"A9",x"FF",x"8D",x"03",x"D3",x"A9",x"BB",x"8D",x"04",x"D1",x"A9",x"F3",x"8D",x"04",x"D2",x"A9",x"8B",x"8D",x"04",x"D3",x"A9",x"55",x"8D",x"05",x"D1",x"A9",x"EC",x"8D",x"05",x"D2",x"A9",x"85",x"8D",x"05",x"D3",x"A9",x"D1",x"8D",x"06",x"D1",x"A9",x"E0",x"8D",x"06",x"D2",x"A9",x"79",x"8D",x"06",x"D3",x"A9",x"AE",x"8D",x"07",x"D1",x"A9",x"5F",x"8D",x"07",x"D2",x"A9",x"C7",x"8D",x"07",x"D3",x"A9",x"9B",x"8D",x"08",x"D1",x"A9",x"47",x"8D",x"08",x"D2",x"A9",x"81",x"8D",x"08",x"D3",x"A9",x"87",x"8D",x"09",x"D1",x"A9",x"37",x"8D",x"09",x"D2",x"A9",x"00",x"8D",x"09",x"D3",x"A9",x"DD",x"8D",x"0A",x"D1",x"A9",x"39",x"8D",x"0A",x"D2",x"A9",x"78",x"8D",x"0A",x"D3",x"A9",x"B5",x"8D",x"0B",x"D1",x"8D",x"0B",x"D2",x"8D",x"0B",x"D3",x"A9",x"B8",x"8D",x"0C",x"D1",x"8D",x"0C",x"D2",x"8D",x"0C",x"D3",x"A9",x"0B",x"8D",x"0D",x"D1",x"A9",x"4F",x"8D",x"0D",x"D2",x"A9",x"CA",x"8D",x"0D",x"D3",x"A9",x"AA",x"8D",x"0E",x"D1",x"A9",x"D9",x"8D",x"0E",x"D2",x"A9",x"FE",x"8D",x"0E",x"D3",x"A9",x"8B",x"8D",x"0F",x"D1",x"8D",x"0F",x"D2",x"8D",x"0F",x"D3",x"A2",x"10",x"8A",x"4A",x"4A",x"4A",x"29",x"0E",x"9D",x"00",x"D1",x"8A",x"4A",x"29",x"0E",x"9D",x"00",x"D2",x"8A",x"0A",x"0A",x"29",x"0C",x"9D",x"00",x"D3",x"E8",x"D0",x"E5",x"60",x"A9",x"01",x"0C",x"30",x"D0",x"A9",x"20",x"8D",x"00",x"04",x"8D",x"02",x"04",x"A9",x"00",x"8D",x"01",x"04",x"8D",x"03",x"04",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"00",x"8D",x"05",x"D7",x"A9",x"00",x"8D",x"06",x"D7",x"A9",x"93",x"8D",x"01",x"D7",x"A9",x"FD",x"8D",x"00",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"8D",x"05",x"D7",x"A9",x"00",x"8D",x"06",x"D7",x"A9",x"94",x"8D",x"01",x"D7",x"A9",x"1E",x"8D",x"00",x"D7",x"A9",x"00",x"8D",x"05",x"D7",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"08",x"8D",x"01",x"CE",x"A2",x"00",x"A0",x"00",x"8A",x"99",x"00",x"04",x"09",x"08",x"99",x"50",x"04",x"8A",x"09",x"10",x"99",x"A0",x"04",x"8A",x"09",x"18",x"99",x"F0",x"04",x"8A",x"09",x"20",x"99",x"40",x"05",x"8A",x"09",x"28",x"99",x"90",x"05",x"8A",x"09",x"30",x"99",x"E0",x"05",x"8A",x"09",x"38",x"99",x"30",x"06",x"C8",x"C8",x"E8",x"E0",x"08",x"D0",x"CC",x"A2",x"00",x"A9",x"01",x"9D",x"01",x"04",x"9D",x"51",x"04",x"9D",x"A1",x"04",x"9D",x"F1",x"04",x"9D",x"41",x"05",x"9D",x"91",x"05",x"9D",x"E1",x"05",x"9D",x"31",x"06",x"E8",x"E8",x"E0",x"10",x"D0",x"E2",x"A9",x"FF",x"8D",x"4E",x"04",x"8D",x"4F",x"04",x"8D",x"9E",x"04",x"8D",x"9F",x"04",x"8D",x"EE",x"04",x"8D",x"EF",x"04",x"8D",x"3E",x"05",x"8D",x"3F",x"05",x"8D",x"8E",x"05",x"8D",x"8F",x"05",x"8D",x"DE",x"05",x"8D",x"DF",x"05",x"8D",x"2E",x"06",x"8D",x"2F",x"06",x"8D",x"7E",x"06",x"8D",x"7F",x"06",x"60",x"04",x"CC",x"07",x"00",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"07",x"D0",x"07",x"01",x"00",x"00",x"00",x"D8",x"80",x"00",x"00",x"03",x"00",x"10",x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00",x"10",x"04",x"9C",x"0F",x"00",x"C0",x"00",x"00",x"00",x"86",x"0B",x"84",x"0C",x"A9",x"00",x"85",x"0D",x"A9",x"04",x"85",x"0E",x"AE",x"01",x"CE",x"E0",x"19",x"D0",x"05",x"A2",x"08",x"8E",x"01",x"CE",x"E0",x"00",x"F0",x"22",x"18",x"A5",x"0D",x"69",x"50",x"85",x"0D",x"A5",x"0E",x"69",x"00",x"85",x"0E",x"C9",x"0B",x"90",x"0E",x"A5",x"0D",x"C9",x"D0",x"90",x"08",x"A9",x"80",x"85",x"0D",x"A9",x"06",x"85",x"0E",x"CA",x"D0",x"DA",x"A0",x"00",x"A9",x"20",x"91",x"0D",x"C8",x"A9",x"00",x"91",x"0D",x"C8",x"C0",x"50",x"D0",x"F2",x"DB",x"A0",x"00",x"A3",x"00",x"B1",x"0B",x"F0",x"13",x"C9",x"40",x"90",x"02",x"29",x"1F",x"92",x"0D",x"1B",x"48",x"A9",x"00",x"92",x"0D",x"68",x"C8",x"1B",x"D0",x"E9",x"EE",x"01",x"CE",x"FB",x"60",x"86",x"0B",x"84",x"0C",x"A9",x"04",x"8D",x"0D",x"BF",x"A9",x"05",x"8D",x"0E",x"BF",x"20",x"77",x"94",x"CE",x"01",x"CE",x"60",x"6B",x"4A",x"4A",x"4A",x"4A",x"20",x"B8",x"94",x"6B",x"29",x"0F",x"AA",x"B1",x"0D",x"C9",x"24",x"F0",x"07",x"C8",x"C8",x"C0",x"50",x"D0",x"F4",x"60",x"8A",x"09",x"30",x"C9",x"3A",x"90",x"02",x"E9",x"39",x"91",x"0D",x"C8",x"C8",x"60",x"AD",x"F1",x"D6",x"10",x"0C",x"A2",x"56",x"A0",x"9A",x"20",x"29",x"94",x"AD",x"F1",x"D6",x"30",x"FB",x"A9",x"82",x"8D",x"80",x"D6",x"A2",x"00",x"8A",x"9D",x"00",x"08",x"E8",x"D0",x"FA",x"A9",x"00",x"8D",x"54",x"D0",x"A9",x"28",x"8D",x"40",x"D0",x"A9",x"00",x"8D",x"41",x"D0",x"20",x"76",x"8B",x"20",x"B8",x"8B",x"8D",x"7F",x"D6",x"8D",x"05",x"D7",x"A9",x"FF",x"8D",x"06",x"D7",x"8E",x"34",x"95",x"8C",x"35",x"95",x"9C",x"36",x"95",x"A9",x"95",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"31",x"8D",x"00",x"D7",x"60",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"BC",x"0F",x"00",x"00",x"A9",x"00",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"AA",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"60",x"B0",x"06",x"A9",x"00",x"8D",x"2F",x"D0",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"60",x"A9",x"FF",x"8D",x"03",x"DC",x"A9",x"00",x"8D",x"02",x"DC",x"A9",x"FE",x"8D",x"01",x"DC",x"A9",x"20",x"AE",x"00",x"DC",x"E0",x"7F",x"D0",x"02",x"A9",x"31",x"E0",x"EF",x"D0",x"02",x"A9",x"39",x"E0",x"F7",x"D0",x"02",x"A9",x"37",x"E0",x"FB",x"D0",x"02",x"A9",x"35",x"E0",x"FD",x"D0",x"02",x"A9",x"33",x"A2",x"F7",x"8E",x"01",x"DC",x"AE",x"00",x"DC",x"E0",x"7F",x"D0",x"02",x"A9",x"32",x"E0",x"EF",x"D0",x"02",x"A9",x"30",x"E0",x"F7",x"D0",x"02",x"A9",x"38",x"E0",x"FB",x"D0",x"02",x"A9",x"36",x"E0",x"FD",x"D0",x"02",x"A9",x"34",x"A2",x"05",x"C9",x"20",x"F0",x"04",x"9D",x"D7",x"9B",x"E8",x"A9",x"2E",x"9D",x"D7",x"9B",x"E8",x"A9",x"52",x"9D",x"D7",x"9B",x"E8",x"A9",x"4F",x"9D",x"D7",x"9B",x"E8",x"A9",x"4D",x"9D",x"D7",x"9B",x"60",x"AD",x"F1",x"D6",x"29",x"01",x"D0",x"01",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"A9",x"FF",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"A9",x"80",x"A2",x"8D",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"AD",x"E1",x"D6",x"4A",x"29",x"02",x"09",x"01",x"8D",x"E1",x"D6",x"60",x"AD",x"F1",x"D6",x"29",x"01",x"D0",x"01",x"60",x"AD",x"E1",x"D6",x"29",x"20",x"D0",x"01",x"60",x"AD",x"E1",x"D6",x"29",x"04",x"4A",x"09",x"01",x"8D",x"E1",x"D6",x"A2",x"09",x"BD",x"0E",x"68",x"DD",x"AC",x"96",x"D3",x"54",x"00",x"CA",x"10",x"F4",x"AD",x"2B",x"68",x"C9",x"41",x"D3",x"49",x"00",x"A9",x"2A",x"8D",x"E2",x"D6",x"A9",x"00",x"8D",x"E3",x"D6",x"A2",x"14",x"BD",x"02",x"68",x"9D",x"00",x"68",x"CA",x"10",x"F7",x"A2",x"05",x"BD",x"08",x"68",x"9D",x"00",x"68",x"A9",x"40",x"9D",x"06",x"68",x"9D",x"16",x"68",x"CA",x"10",x"EF",x"A9",x"02",x"8D",x"15",x"68",x"A2",x"03",x"BD",x"28",x"68",x"9D",x"1C",x"68",x"CA",x"10",x"F7",x"A2",x"09",x"BD",x"18",x"68",x"9D",x"20",x"68",x"CA",x"10",x"F7",x"A9",x"01",x"8D",x"E4",x"D6",x"AD",x"10",x"68",x"C9",x"45",x"D0",x"1F",x"AD",x"19",x"68",x"C9",x"11",x"D0",x"18",x"AD",x"26",x"68",x"C9",x"11",x"D0",x"11",x"AD",x"27",x"68",x"C9",x"9F",x"D0",x"0A",x"AD",x"2C",x"68",x"C9",x"A9",x"D0",x"03",x"20",x"2C",x"68",x"60",x"08",x"06",x"00",x"01",x"08",x"00",x"06",x"04",x"00",x"01",x"C9",x"0A",x"B0",x"03",x"09",x"30",x"60",x"38",x"E9",x"09",x"60",x"08",x"DB",x"5A",x"DA",x"48",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"82",x"06",x"68",x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"80",x"06",x"AD",x"F9",x"BC",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"84",x"06",x"AD",x"F9",x"BC",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"86",x"06",x"AD",x"84",x"D6",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"8A",x"06",x"AD",x"84",x"D6",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"8C",x"06",x"AD",x"83",x"D6",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"8E",x"06",x"AD",x"83",x"D6",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"90",x"06",x"AD",x"82",x"D6",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"92",x"06",x"AD",x"82",x"D6",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"94",x"06",x"AD",x"81",x"D6",x"4A",x"4A",x"4A",x"4A",x"20",x"B6",x"96",x"8D",x"96",x"06",x"AD",x"81",x"D6",x"29",x"0F",x"20",x"B6",x"96",x"8D",x"98",x"06",x"AD",x"F1",x"D6",x"AE",x"F0",x"D6",x"CD",x"F1",x"D6",x"D0",x"0B",x"EC",x"F0",x"D6",x"D0",x"06",x"EE",x"20",x"D0",x"4C",x"58",x"97",x"A2",x"00",x"A0",x"00",x"A3",x"F0",x"E8",x"D0",x"FD",x"C8",x"D0",x"FA",x"1B",x"D0",x"F7",x"68",x"FA",x"7A",x"FB",x"28",x"60",x"43",x"36",x"35",x"47",x"53",x"20",x"4B",x"49",x"43",x"4B",x"53",x"54",x"41",x"52",x"54",x"20",x"56",x"30",x"30",x"2E",x"30",x"33",x"00",x"52",x"4F",x"4D",x"20",x"43",x"48",x"45",x"43",x"4B",x"53",x"55",x"4D",x"20",x"4F",x"4B",x"20",x"2D",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"00",x"52",x"4F",x"4D",x"20",x"43",x"48",x"45",x"43",x"4B",x"53",x"55",x"4D",x"20",x"46",x"41",x"49",x"4C",x"20",x"2D",x"20",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"52",x"4F",x"4D",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4C",x"4F",x"41",x"44",x"20",x"43",x"48",x"41",x"52",x"52",x"4F",x"4D",x"2E",x"47",x"36",x"35",x"00",x"4C",x"4F",x"41",x"44",x"45",x"44",x"20",x"43",x"48",x"41",x"52",x"52",x"4F",x"4D",x"2E",x"47",x"36",x"35",x"20",x"28",x"24",x"24",x"24",x"24",x"20",x"50",x"41",x"47",x"45",x"53",x"29",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"2E",x"2E",x"2E",x"00",x"46",x"4F",x"55",x"4E",x"44",x"20",x"41",x"4E",x"44",x"20",x"52",x"45",x"53",x"45",x"54",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"00",x"45",x"52",x"52",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"20",x"43",x"41",x"52",x"44",x"00",x"42",x"41",x"44",x"20",x"4D",x"42",x"52",x"20",x"4F",x"52",x"20",x"44",x"4F",x"53",x"20",x"42",x"4F",x"4F",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"2E",x"00",x"52",x"45",x"41",x"44",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"54",x"41",x"42",x"4C",x"45",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"00",x"46",x"4F",x"55",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"20",x"3D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"20",x"24",x"24",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"53",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"24",x"24",x"20",x"42",x"59",x"54",x"45",x"53",x"2C",x"20",x"49",x"20",x"53",x"45",x"45",x"20",x"24",x"24",x"20",x"42",x"59",x"54",x"45",x"53",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4F",x"50",x"45",x"4E",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"20",x"46",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"00",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"2E",x"2E",x"00",x"52",x"4F",x"4D",x"20",x"54",x"4F",x"4F",x"20",x"4C",x"4F",x"4E",x"47",x"3A",x"20",x"28",x"52",x"45",x"41",x"44",x"20",x"24",x"24",x"24",x"24",x"20",x"50",x"41",x"47",x"45",x"53",x"29",x"00",x"52",x"4F",x"4D",x"20",x"54",x"4F",x"4F",x"20",x"53",x"48",x"4F",x"52",x"54",x"3A",x"20",x"28",x"52",x"45",x"41",x"44",x"20",x"24",x"24",x"24",x"24",x"20",x"50",x"41",x"47",x"45",x"53",x"29",x"00",x"20",x"4E",x"45",x"58",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"3D",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"4E",x"45",x"58",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"3D",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"43",x"41",x"4E",x"4E",x"4F",x"54",x"20",x"46",x"49",x"4E",x"44",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"2D",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"20",x"24",x"24",x"29",x"00",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"40",x"20",x"49",x"4E",x"54",x"45",x"52",x"4E",x"41",x"4C",x"20",x"46",x"30",x"31",x"31",x"20",x"44",x"52",x"49",x"56",x"45",x"00",x"46",x"41",x"49",x"4C",x"3A",x"20",x"43",x"36",x"34",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"49",x"53",x"20",x"4E",x"4F",x"54",x"20",x"38",x"31",x"39",x"32",x"30",x"30",x"20",x"42",x"59",x"54",x"45",x"53",x"20",x"4C",x"4F",x"4E",x"47",x"00",x"46",x"41",x"49",x"4C",x"3A",x"20",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"49",x"53",x"20",x"46",x"52",x"41",x"47",x"4D",x"45",x"4E",x"54",x"45",x"44",x"3A",x"20",x"44",x"45",x"46",x"52",x"41",x"47",x"20",x"49",x"54",x"00",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"20",x"53",x"55",x"43",x"43",x"45",x"53",x"53",x"46",x"55",x"4C",x"4C",x"59",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"00",x"52",x"45",x"4C",x"45",x"41",x"53",x"45",x"20",x"53",x"57",x"31",x"35",x"20",x"54",x"4F",x"20",x"43",x"4F",x"4E",x"54",x"49",x"4E",x"55",x"45",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"2E",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"46",x"49",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"43",x"36",x"35",x"47",x"53",x"58",x"58",x"58",x"52",x"4F",x"4D",x"00",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"4B",x"49",x"43",x"4B",x"55",x"50",x"2E",x"47",x"36",x"35",x"20",x"49",x"4E",x"54",x"4F",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"00",x"4E",x"4F",x"20",x"4B",x"49",x"43",x"4B",x"55",x"50",x"2E",x"47",x"36",x"35",x"20",x"54",x"4F",x"20",x"4C",x"4F",x"41",x"44",x"20",x"28",x"4F",x"52",x"20",x"42",x"52",x"4F",x"4B",x"45",x"4E",x"29",x"00",x"4B",x"49",x"43",x"4B",x"55",x"50",x"20",x"4C",x"4F",x"41",x"44",x"45",x"44",x"20",x"54",x"4F",x"20",x"30",x"30",x"30",x"30",x"34",x"30",x"30",x"30",x"20",x"2D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"52",x"55",x"4E",x"4E",x"49",x"4E",x"47",x"20",x"4B",x"49",x"43",x"4B",x"45",x"44",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"00",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"20",x"56",x"49",x"41",x"20",x"45",x"54",x"48",x"45",x"52",x"4B",x"49",x"43",x"4B",x"3A",x"20",x"55",x"44",x"50",x"20",x"50",x"4F",x"52",x"54",x"20",x"34",x"35",x"31",x"31",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"4E",x"45",x"58",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"20",x"4F",x"46",x"20",x"46",x"49",x"4C",x"45",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4C",x"4F",x"41",x"44",x"20",x"42",x"4F",x"4F",x"54",x"4C",x"4F",x"47",x"4F",x"2E",x"47",x"36",x"35",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"24",x"24",x"29",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"43",x"48",x"44",x"49",x"52",x"20",x"54",x"4F",x"20",x"2F",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"24",x"24",x"29",x"00",x"47",x"49",x"54",x"20",x"43",x"4F",x"4D",x"4D",x"49",x"54",x"3A",x"20",x"46",x"41",x"39",x"45",x"42",x"34",x"38",x"33",x"43",x"41",x"46",x"35",x"46",x"38",x"41",x"2A",x"2B",x"44",x"49",x"52",x"54",x"59",x"00",x"00",x"43",x"48",x"41",x"52",x"52",x"4F",x"4D",x"2E",x"47",x"36",x"35",x"00",x"43",x"36",x"35",x"47",x"53",x"2E",x"52",x"4F",x"4D",x"00",x"00",x"43",x"36",x"35",x"47",x"53",x"2E",x"44",x"38",x"31",x"00",x"4B",x"49",x"43",x"4B",x"55",x"50",x"2E",x"47",x"36",x"35",x"00",x"42",x"4F",x"4F",x"54",x"4C",x"4F",x"47",x"4F",x"2E",x"47",x"36",x"35",x"00",x"BA",x"8E",x"5A",x"CE",x"A9",x"93",x"20",x"D2",x"FF",x"38",x"20",x"DC",x"C6",x"78",x"20",x"AC",x"C6",x"4F",x"50",x"45",x"4E",x"49",x"4E",x"47",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"2E",x"2E",x"2E",x"0D",x"00",x"20",x"5E",x"C5",x"B0",x"03",x"4C",x"24",x"C0",x"20",x"AC",x"C6",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"54",x"41",x"42",x"4C",x"45",x"2E",x"2E",x"2E",x"0D",x"00",x"20",x"EC",x"C5",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"DB",x"02",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"D3",x"02",x"A0",x"00",x"AB",x"C9",x"DF",x"9C",x"0B",x"CE",x"AB",x"C8",x"DF",x"9C",x"0A",x"CE",x"AB",x"C7",x"DF",x"9C",x"09",x"CE",x"AB",x"C6",x"DF",x"9C",x"08",x"CE",x"A2",x"03",x"BD",x"08",x"CE",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"20",x"77",x"C6",x"20",x"FA",x"C5",x"93",x"90",x"02",x"20",x"AC",x"C6",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"2E",x"2E",x"2E",x"0D",x"00",x"AD",x"FE",x"DF",x"C9",x"55",x"D3",x"83",x"02",x"AD",x"FF",x"DF",x"C9",x"AA",x"D3",x"7B",x"02",x"AD",x"11",x"DE",x"D3",x"75",x"02",x"A2",x"03",x"BD",x"0E",x"DE",x"9D",x"10",x"CE",x"9D",x"0C",x"CE",x"BD",x"2C",x"DE",x"9D",x"14",x"CE",x"CA",x"10",x"EE",x"A9",x"00",x"8D",x"12",x"CE",x"8D",x"13",x"CE",x"8D",x"0E",x"CE",x"8D",x"0F",x"CE",x"AC",x"10",x"DE",x"F0",x"18",x"A2",x"00",x"18",x"08",x"28",x"BD",x"10",x"CE",x"7D",x"24",x"DE",x"9D",x"10",x"CE",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"88",x"D0",x"E8",x"38",x"A2",x"03",x"BD",x"20",x"DE",x"FD",x"10",x"CE",x"9D",x"1C",x"CE",x"9D",x"20",x"CE",x"CA",x"10",x"F1",x"AD",x"0D",x"DE",x"8D",x"24",x"CE",x"A8",x"29",x"FE",x"F0",x"14",x"A2",x"03",x"18",x"BD",x"20",x"CE",x"6A",x"9D",x"20",x"CE",x"CA",x"10",x"F6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"AD",x"23",x"CE",x"0D",x"22",x"CE",x"F3",x"FC",x"01",x"A2",x"03",x"BD",x"2C",x"DE",x"9D",x"18",x"CE",x"9D",x"4A",x"CE",x"CA",x"10",x"F4",x"20",x"AC",x"C6",x"53",x"45",x"41",x"52",x"43",x"48",x"49",x"4E",x"47",x"20",x"44",x"49",x"52",x"45",x"43",x"54",x"4F",x"52",x"59",x"2E",x"2E",x"2E",x"0D",x"00",x"A9",x"00",x"8D",x"8B",x"D6",x"20",x"78",x"C3",x"20",x"87",x"C3",x"93",x"B0",x"01",x"EA",x"20",x"9C",x"C3",x"93",x"79",x"01",x"A2",x"00",x"AD",x"31",x"CE",x"20",x"6D",x"C3",x"C9",x"44",x"D0",x"ED",x"AD",x"32",x"CE",x"20",x"6D",x"C3",x"C9",x"38",x"D0",x"E3",x"AD",x"33",x"CE",x"20",x"6D",x"C3",x"C9",x"31",x"D0",x"D9",x"20",x"AC",x"C6",x"4D",x"4F",x"55",x"4E",x"54",x"20",x"00",x"20",x"F3",x"C5",x"A2",x"00",x"BD",x"29",x"CE",x"DA",x"20",x"D2",x"FF",x"FA",x"E8",x"E0",x"08",x"D0",x"F3",x"20",x"AC",x"C6",x"3F",x"20",x"00",x"20",x"F3",x"C5",x"58",x"20",x"E4",x"FF",x"C9",x"00",x"F0",x"F9",x"48",x"A9",x"0D",x"20",x"D2",x"FF",x"78",x"20",x"EC",x"C5",x"68",x"C9",x"59",x"D0",x"9D",x"20",x"EB",x"C3",x"20",x"EE",x"C4",x"20",x"77",x"C6",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"8C",x"D6",x"CA",x"10",x"F7",x"20",x"EB",x"C3",x"A2",x"03",x"BD",x"4A",x"CE",x"9D",x"4F",x"CE",x"CA",x"10",x"F7",x"A9",x"00",x"8D",x"55",x"CE",x"8D",x"56",x"CE",x"A9",x"40",x"8D",x"53",x"CE",x"A9",x"06",x"8D",x"54",x"CE",x"AB",x"24",x"CE",x"6B",x"29",x"01",x"D0",x"0C",x"6B",x"4A",x"4B",x"4E",x"54",x"CE",x"6E",x"53",x"CE",x"4C",x"06",x"C2",x"A2",x"03",x"BD",x"4F",x"CE",x"DD",x"4A",x"CE",x"D3",x"81",x"00",x"CA",x"10",x"F4",x"EE",x"55",x"CE",x"D0",x"03",x"EE",x"56",x"CE",x"18",x"AD",x"4F",x"CE",x"69",x"01",x"8D",x"4F",x"CE",x"AD",x"50",x"CE",x"69",x"00",x"8D",x"50",x"CE",x"AD",x"51",x"CE",x"69",x"00",x"8D",x"51",x"CE",x"AD",x"52",x"CE",x"69",x"00",x"8D",x"52",x"CE",x"20",x"38",x"C4",x"B0",x"C4",x"AD",x"53",x"CE",x"CD",x"55",x"CE",x"D0",x"25",x"AD",x"54",x"CE",x"CD",x"56",x"CE",x"D0",x"1D",x"A9",x"07",x"8D",x"8B",x"D6",x"18",x"20",x"DC",x"C6",x"20",x"AC",x"C6",x"44",x"49",x"53",x"4B",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"2E",x"44",x"38",x"31",x"20",x"46",x"49",x"4C",x"45",x"20",x"48",x"41",x"53",x"20",x"57",x"52",x"4F",x"4E",x"47",x"20",x"4C",x"45",x"4E",x"47",x"54",x"48",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"54",x"48",x"41",x"54",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"20",x"49",x"53",x"20",x"46",x"52",x"41",x"47",x"4D",x"45",x"4E",x"54",x"45",x"44",x"2E",x"0D",x"44",x"45",x"2D",x"46",x"52",x"41",x"47",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"20",x"42",x"45",x"46",x"4F",x"52",x"45",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"49",x"4E",x"47",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"4E",x"4F",x"20",x"4D",x"4F",x"52",x"45",x"20",x"44",x"49",x"53",x"4B",x"20",x"49",x"4D",x"41",x"47",x"45",x"53",x"2E",x"20",x"44",x"52",x"49",x"56",x"45",x"20",x"4D",x"41",x"52",x"4B",x"45",x"44",x"20",x"45",x"4D",x"50",x"54",x"59",x"2E",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"53",x"44",x"2D",x"43",x"41",x"52",x"44",x"20",x"45",x"52",x"52",x"4F",x"52",x"0D",x"00",x"4C",x"EF",x"C6",x"20",x"AC",x"C6",x"49",x"4E",x"56",x"41",x"4C",x"49",x"44",x"20",x"4F",x"52",x"20",x"55",x"4E",x"53",x"55",x"50",x"50",x"4F",x"52",x"54",x"45",x"44",x"20",x"46",x"49",x"4C",x"45",x"20",x"53",x"59",x"53",x"54",x"45",x"4D",x"2E",x"0D",x"28",x"53",x"48",x"4F",x"55",x"4C",x"44",x"20",x"42",x"45",x"20",x"46",x"41",x"54",x"33",x"32",x"29",x"0D",x"00",x"4C",x"EF",x"C6",x"C9",x"60",x"90",x"06",x"C9",x"7A",x"B0",x"02",x"29",x"5F",x"60",x"A2",x"00",x"BD",x"18",x"CE",x"9D",x"25",x"CE",x"E8",x"E0",x"04",x"D0",x"F5",x"38",x"60",x"A2",x"00",x"BD",x"25",x"CE",x"9D",x"4A",x"CE",x"E8",x"E0",x"04",x"D0",x"F5",x"A9",x"00",x"8D",x"49",x"CE",x"4C",x"05",x"C4",x"AD",x"49",x"CE",x"C9",x"10",x"90",x"0B",x"A9",x"00",x"8D",x"49",x"CE",x"20",x"16",x"C4",x"B0",x"01",x"60",x"A0",x"00",x"AD",x"49",x"CE",x"29",x"08",x"D0",x"1A",x"AD",x"49",x"CE",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DE",x"99",x"29",x"CE",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CE",x"38",x"60",x"AD",x"49",x"CE",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"BD",x"00",x"DF",x"99",x"29",x"CE",x"E8",x"C8",x"C0",x"20",x"D0",x"F4",x"EE",x"49",x"CE",x"38",x"60",x"AD",x"3D",x"CE",x"8D",x"4C",x"CE",x"AD",x"3E",x"CE",x"8D",x"4D",x"CE",x"AD",x"43",x"CE",x"8D",x"4A",x"CE",x"AD",x"44",x"CE",x"8D",x"4B",x"CE",x"38",x"60",x"A9",x"00",x"8D",x"4E",x"CE",x"20",x"EE",x"C4",x"B0",x"01",x"60",x"20",x"77",x"C6",x"4C",x"FA",x"C5",x"20",x"43",x"C6",x"EE",x"4E",x"CE",x"AD",x"4E",x"CE",x"CD",x"24",x"CE",x"D0",x"11",x"A9",x"00",x"8D",x"4E",x"CE",x"20",x"38",x"C4",x"B0",x"01",x"60",x"20",x"EE",x"C4",x"20",x"77",x"C6",x"4C",x"FA",x"C5",x"A2",x"00",x"BD",x"4A",x"CE",x"9D",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F5",x"A0",x"07",x"18",x"6E",x"84",x"D6",x"6E",x"83",x"D6",x"6E",x"82",x"D6",x"6E",x"81",x"D6",x"88",x"D0",x"F0",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CE",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"0C",x"CE",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"20",x"77",x"C6",x"20",x"FA",x"C5",x"90",x"63",x"AD",x"4A",x"CE",x"0A",x"0A",x"AA",x"A0",x"00",x"AD",x"4A",x"CE",x"29",x"40",x"D0",x"0E",x"BD",x"00",x"DE",x"99",x"4A",x"CE",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"80",x"0C",x"BD",x"00",x"DF",x"99",x"4A",x"CE",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"AD",x"4D",x"CE",x"29",x"0F",x"8D",x"4D",x"CE",x"AD",x"4D",x"CE",x"0D",x"4C",x"CE",x"0D",x"4B",x"CE",x"0D",x"4A",x"CE",x"C9",x"00",x"F0",x"22",x"AD",x"4D",x"CE",x"C9",x"0F",x"D0",x"19",x"AD",x"4C",x"CE",x"C9",x"FF",x"D0",x"12",x"AD",x"4B",x"CE",x"C9",x"FF",x"D0",x"0B",x"AD",x"4A",x"CE",x"C9",x"FF",x"F0",x"06",x"C9",x"F7",x"F0",x"02",x"38",x"60",x"18",x"60",x"A2",x"03",x"BD",x"4A",x"CE",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A2",x"03",x"38",x"08",x"28",x"BD",x"81",x"D6",x"FD",x"14",x"CE",x"9D",x"81",x"D6",x"08",x"CA",x"10",x"F2",x"28",x"AD",x"24",x"CE",x"A8",x"29",x"FE",x"F0",x"14",x"18",x"2E",x"81",x"D6",x"2E",x"82",x"D6",x"2E",x"83",x"D6",x"2E",x"84",x"D6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"A2",x"00",x"BD",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"10",x"CE",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"7D",x"08",x"CE",x"9D",x"81",x"D6",x"08",x"E8",x"E0",x"04",x"D0",x"F0",x"28",x"38",x"60",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"4C",x"FA",x"C5",x"A9",x"42",x"8D",x"80",x"D6",x"A9",x"00",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F9",x"60",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F9",x"60",x"20",x"AF",x"C5",x"20",x"EC",x"C5",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"AD",x"80",x"D6",x"20",x"D0",x"C5",x"B0",x"03",x"D0",x"F6",x"60",x"38",x"60",x"20",x"C2",x"C5",x"EE",x"57",x"CE",x"D0",x"FB",x"EE",x"58",x"CE",x"D0",x"F6",x"EE",x"59",x"CE",x"D0",x"F1",x"60",x"A9",x"00",x"8D",x"57",x"CE",x"8D",x"58",x"CE",x"A9",x"E0",x"8D",x"59",x"CE",x"60",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"13",x"EE",x"57",x"CE",x"D0",x"0C",x"EE",x"58",x"CE",x"D0",x"07",x"EE",x"59",x"CE",x"D0",x"02",x"A9",x"00",x"18",x"60",x"38",x"60",x"A9",x"81",x"8D",x"80",x"D6",x"38",x"60",x"A9",x"82",x"8D",x"80",x"D6",x"38",x"60",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"40",x"4C",x"16",x"C6",x"EE",x"20",x"D0",x"A2",x"F0",x"A0",x"00",x"A3",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"E8",x"D0",x"F7",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"C2",x"C5",x"20",x"D0",x"C5",x"B0",x"05",x"D0",x"F9",x"4C",x"3B",x"C6",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"EF",x"AD",x"88",x"D6",x"AD",x"89",x"D6",x"C9",x"02",x"D0",x"CB",x"38",x"60",x"20",x"6F",x"C5",x"4C",x"16",x"C6",x"18",x"60",x"AD",x"80",x"D6",x"29",x"10",x"D0",x"1A",x"AD",x"82",x"D6",x"18",x"69",x"02",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"69",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"69",x"00",x"8D",x"84",x"D6",x"60",x"EE",x"81",x"D6",x"90",x"0D",x"EE",x"82",x"D6",x"90",x"08",x"EE",x"83",x"D6",x"90",x"03",x"EE",x"84",x"D6",x"60",x"AD",x"80",x"D6",x"29",x"10",x"F0",x"01",x"60",x"AD",x"83",x"D6",x"8D",x"84",x"D6",x"AD",x"82",x"D6",x"8D",x"83",x"D6",x"AD",x"81",x"D6",x"8D",x"82",x"D6",x"A9",x"00",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"0A",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"2A",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"2A",x"8D",x"84",x"D6",x"60",x"20",x"F3",x"C5",x"58",x"68",x"8D",x"BB",x"C6",x"68",x"8D",x"BC",x"C6",x"A2",x"01",x"BD",x"FF",x"FF",x"F0",x"06",x"20",x"D2",x"FF",x"E8",x"D0",x"F5",x"38",x"8A",x"6D",x"BB",x"C6",x"8D",x"DA",x"C6",x"A9",x"00",x"6D",x"BC",x"C6",x"8D",x"DB",x"C6",x"78",x"20",x"EC",x"C5",x"4C",x"FF",x"FF",x"B0",x"06",x"A9",x"00",x"8D",x"2F",x"D0",x"60",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"60",x"20",x"F3",x"C5",x"18",x"20",x"DC",x"C6",x"AE",x"5A",x"CE",x"9A",x"A9",x"00",x"58",x"18",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"CF",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"A9",x"FF",x"A2",x"0F",x"A0",x"00",x"A3",x"00",x"5C",x"EA",x"A9",x"80",x"A2",x"8D",x"A0",x"00",x"A3",x"00",x"5C",x"EA",x"AD",x"E1",x"D6",x"4A",x"29",x"02",x"09",x"01",x"8D",x"E1",x"D6",x"AD",x"E1",x"D6",x"29",x"20",x"F0",x"F9",x"AD",x"E1",x"D6",x"29",x"04",x"4A",x"09",x"01",x"8D",x"E1",x"D6",x"A2",x"09",x"BD",x"0E",x"68",x"DD",x"CB",x"CF",x"D0",x"52",x"CA",x"10",x"F5",x"AD",x"2B",x"68",x"C9",x"41",x"D0",x"48",x"A9",x"2A",x"8D",x"E2",x"D6",x"A9",x"00",x"8D",x"E3",x"D6",x"A2",x"14",x"BD",x"02",x"68",x"9D",x"00",x"68",x"CA",x"10",x"F7",x"A2",x"05",x"BD",x"08",x"68",x"9D",x"00",x"68",x"A9",x"40",x"9D",x"06",x"68",x"9D",x"16",x"68",x"CA",x"10",x"EF",x"A9",x"02",x"8D",x"15",x"68",x"A2",x"03",x"BD",x"28",x"68",x"9D",x"1C",x"68",x"CA",x"10",x"F7",x"A2",x"09",x"BD",x"18",x"68",x"9D",x"20",x"68",x"CA",x"10",x"F7",x"A9",x"01",x"8D",x"E4",x"D6",x"AD",x"10",x"68",x"C9",x"45",x"D0",x"8B",x"AD",x"19",x"68",x"C9",x"11",x"D0",x"84",x"AD",x"26",x"68",x"C9",x"11",x"D3",x"7D",x"FF",x"AD",x"27",x"68",x"C9",x"9E",x"D3",x"75",x"FF",x"AD",x"2C",x"68",x"C9",x"A9",x"D3",x"6D",x"FF",x"20",x"2C",x"68",x"4C",x"31",x"CF",x"08",x"06",x"00",x"01",x"08",x"00",x"06",x"04",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"56",x"65",x"6E",x"65",x"7A",x"75",x"61",x"6C",x"65",x"6E",x"20",x"63",x"61",x"73",x"61",x"62",x"61",x"20",x"6D",x"65",x"6C",x"6F",x"6E",x"20",x"70",x"72",x"6F",x"64",x"75",x"63",x"74",x"69",x"6F",x"6E",x"20",x"73",x"74",x"61",x"74",x"69",x"73",x"74",x"69",x"63",x"73",x"20",x"28",x"32",x"30",x"31",x"32",x"2D",x"32",x"30",x"31",x"35",x"29",x"2E",x"74",x"78",x"74",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"46",x"49",x"4C",x"45",x"4E",x"41",x"4D",x"45",x"2E",x"45",x"58",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"56",x"65",x"6E",x"65",x"7A",x"75",x"61",x"6C",x"65",x"6E",x"20",x"63",x"61",x"73",x"61",x"62",x"61",x"20",x"6D",x"65",x"6C",x"6F",x"6E",x"20",x"70",x"72",x"6F",x"64",x"75",x"63",x"74",x"69",x"6F",x"6E",x"20",x"73",x"74",x"61",x"74",x"69",x"73",x"74",x"69",x"63",x"73",x"20",x"28",x"32",x"30",x"30",x"37",x"2D",x"32",x"30",x"31",x"31",x"29",x"2E",x"74",x"78",x"74",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"4F",x"50",x"45",x"52",x"41",x"54",x"49",x"4E",x"47",x"20",x"53",x"59",x"53",x"54",x"45",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F");

begin

--process for read and write operation.
  PROCESS(Clk,cs,ram,address)
  BEGIN
    if(rising_edge(Clk)) then 
      if cs='1' then
        if(we='1') then
          ram(to_integer(unsigned(address))) <= data_i;
        end if;
        data_o <= ram(to_integer(unsigned(address)));
      end if;
    end if;
    if cs='1' then
      data_o <= ram(to_integer(unsigned(address)));
    else
      data_o <= "ZZZZZZZZ";
    end if;
  END PROCESS;

end Behavioral;
