vga/vga.vhd