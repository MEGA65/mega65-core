library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use STD.textio.all;
use work.debugtools.all;
use work.cputypes.all;

entity test_buffereduart is
end entity;

architecture foo of test_buffereduart is

  signal cpuclock : std_logic := '1';
  
  signal cycles : integer := 0;

  type mem_transaction_t is record
    address : unsigned(15 downto 0);
    write_p : std_logic;
    value : unsigned(7 downto 0);     -- either to write, or expected to read
    delay : integer;
  end record mem_transaction_t;

  type mem_job_list_t is array(0 to 2047) of mem_transaction_t;

  signal fastio_addr : unsigned(19 downto 0) := to_unsigned(0,20);
  signal fastio_rdata : unsigned(7 downto 0);
  signal fastio_wdata : unsigned(7 downto 0) := x"00";
  signal fastio_write : std_logic := '0';
  signal fastio_read : std_logic := '0';

  signal buffereduart_cs : std_logic := '1';
  signal uart_irq : std_logic := '1';
  signal reset : std_logic := '1';

  signal buffereduart_rx : std_logic_vector(7 downto 0) := (others => '1');
  signal buffereduart_tx : std_logic_vector(7 downto 0) := (others => '1');
  signal buffereduart_ringindicate : std_logic_vector(7 downto 0) := (others => '1');
  
  signal start_time : integer := 0;
  signal current_time : integer := 0;
  signal dispatch_time : integer := 0;
  
  signal mem_jobs : mem_job_list_t := (
    -- Read $D0E0 status register and wait a while for flags to all update
    ( address => x"D0E0", write_p => '0', value => x"00", delay => 0),
    -- Read $D0E1 status register
    ( address => x"D0E1", write_p => '0', value => x"60", delay => 0),

    -- Enable loopback mode for testing, select uart #7
    -- (which will be connected to UART #0 via the loopback)
    ( address => x"D0E0", write_p => '1', value => x"17", delay => 0),    
    
    -- Set data rate for uart #1 very fast for testing
    ( address => x"D0E4", write_p => '1', value => x"04", delay => 0),
    ( address => x"D0E5", write_p => '1', value => x"00", delay => 0),
    ( address => x"D0E6", write_p => '1', value => x"00", delay => 0),        
    
    -- Enable loopback mode for testing, select uart #0
    ( address => x"D0E0", write_p => '1', value => x"10", delay => 0),    
    
    -- Set data rate for uart #0 very fast for testing
    ( address => x"D0E4", write_p => '1', value => x"04", delay => 0),
    ( address => x"D0E5", write_p => '1', value => x"00", delay => 0),
    ( address => x"D0E6", write_p => '1', value => x"00", delay => 0),

    -- Write a char to uart #0, which should then get received by uart #7
    ( address => x"D0E3", write_p => '1', value => x"12", delay => 2),
    -- Read at the right time to observe that tx_empty is cleared
    ( address => x"D0E1", write_p => '0', value => x"40", delay => 8),
    -- Read at the right time to observe that tx_empty is again asserted
    ( address => x"D0E1", write_p => '0', value => x"60", delay => 0),

    -- Now select uart #7, and see what we can see there
    -- We add a delay of 70 cycles to allow for the RX of the byte to complete
    ( address => x"D0E0", write_p => '1', value => x"17", delay => 70),
    
    -- rx_empty should be clear
    ( address => x"D0E1", write_p => '0', value => x"20", delay => 0),
    -- see if we can read the received byte ok
    ( address => x"D0E2", write_p => '0', value => x"12", delay => 0),
    -- Acknowledge the received byte
    ( address => x"D0E2", write_p => '1', value => x"00", delay => 8),
    -- rx_empty should be asserted again now
    ( address => x"D0E1", write_p => '0', value => x"60", delay => 0),

    -- Now send two more bytes
    ( address => x"D0E0", write_p => '1', value => x"10", delay => 0),    
    ( address => x"D0E3", write_p => '1', value => x"34", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"56", delay => 2),
    ( address => x"D0E0", write_p => '1', value => x"17", delay => 200),
    ( address => x"D0E1", write_p => '0', value => x"20", delay => 0),
    ( address => x"D0E2", write_p => '0', value => x"34", delay => 0),
    ( address => x"D0E2", write_p => '1', value => x"00", delay => 8),
    ( address => x"D0E2", write_p => '0', value => x"56", delay => 0),
    ( address => x"D0E2", write_p => '1', value => x"00", delay => 8),
    ( address => x"D0E1", write_p => '0', value => x"60", delay => 0),

    -- Send lots of bytes, and wait for TX low-water to clear
    ( address => x"D0E0", write_p => '1', value => x"10", delay => 0),    

    ( address => x"D0E3", write_p => '1', value => x"00", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"01", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"02", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"03", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"04", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"05", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"06", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"07", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"08", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"09", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"0f", delay => 2),

    ( address => x"D0E3", write_p => '1', value => x"10", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"11", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"12", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"13", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"14", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"15", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"16", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"17", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"18", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"19", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"1f", delay => 2),

    ( address => x"D0E3", write_p => '1', value => x"20", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"21", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"22", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"23", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"24", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"25", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"26", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"27", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"28", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"29", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"2f", delay => 2),
    
    ( address => x"D0E3", write_p => '1', value => x"30", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"31", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"32", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"33", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"34", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"35", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"36", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"37", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"38", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"39", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"3f", delay => 2),
    
    ( address => x"D0E3", write_p => '1', value => x"40", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"41", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"42", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"43", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"44", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"45", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"46", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"47", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"48", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"49", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"4f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"50", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"51", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"52", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"53", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"54", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"55", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"56", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"57", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"58", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"59", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"5f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"60", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"61", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"62", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"63", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"64", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"65", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"66", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"67", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"68", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"69", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"6f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"70", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"71", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"72", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"73", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"74", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"75", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"76", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"77", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"78", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"79", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"7f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"80", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"81", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"82", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"83", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"84", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"85", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"86", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"87", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"88", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"89", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"8f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"90", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"91", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"92", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"93", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"94", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"95", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"96", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"97", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"98", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"99", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9a", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9b", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9c", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9d", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9e", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"9f", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"a9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"aa", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ab", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ac", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ad", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ae", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"af", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"b9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ba", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"bb", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"bc", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"bd", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"be", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"bf", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"c9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ca", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"cb", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"cc", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"cd", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ce", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"cf", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"d9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"da", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"db", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"dc", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"dd", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"de", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"df", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"e9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ea", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"eb", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ec", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ed", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ee", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ef", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f0", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f1", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f2", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f3", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f4", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f5", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f6", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f7", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f8", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"f9", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"fa", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"fb", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"fc", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"fd", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"fe", delay => 2),
    ( address => x"D0E3", write_p => '1', value => x"ff", delay => 2),

    -- Now select uart #7 again, and read all those bytes out
    -- (and allow enough delay for each to be received
    ( address => x"D0E0", write_p => '1', value => x"17", delay => 0),
    
    
    ( address => x"D0E2", write_p => '0', value => x"00", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"00", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"01", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"01", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"02", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"02", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"03", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"03", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"04", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"04", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"05", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"05", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"06", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"06", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"07", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"07", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"08", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"08", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"09", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"09", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"0f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"0f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"10", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"10", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"11", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"11", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"12", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"12", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"13", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"13", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"14", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"14", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"15", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"15", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"16", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"16", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"17", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"17", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"18", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"18", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"19", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"19", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"1f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"1f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"20", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"20", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"21", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"21", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"22", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"22", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"23", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"23", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"24", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"24", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"25", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"25", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"26", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"26", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"27", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"27", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"28", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"28", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"29", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"29", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"2f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"2f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"30", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"30", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"31", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"31", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"32", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"32", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"33", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"33", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"34", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"34", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"35", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"35", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"36", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"36", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"37", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"37", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"38", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"38", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"39", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"39", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"3f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"3f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"40", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"40", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"41", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"41", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"42", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"42", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"43", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"43", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"44", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"44", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"45", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"45", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"46", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"46", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"47", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"47", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"48", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"48", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"49", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"49", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"4f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"4f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"50", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"50", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"51", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"51", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"52", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"52", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"53", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"53", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"54", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"54", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"55", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"55", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"56", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"56", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"57", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"57", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"58", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"58", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"59", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"59", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"5f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"5f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"60", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"60", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"61", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"61", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"62", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"62", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"63", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"63", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"64", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"64", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"65", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"65", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"66", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"66", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"67", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"67", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"68", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"68", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"69", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"69", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"6f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"6f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"70", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"70", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"71", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"71", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"72", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"72", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"73", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"73", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"74", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"74", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"75", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"75", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"76", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"76", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"77", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"77", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"78", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"78", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"79", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"79", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"7f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"7f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"80", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"80", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"81", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"81", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"82", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"82", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"83", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"83", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"84", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"84", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"85", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"85", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"86", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"86", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"87", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"87", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"88", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"88", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"89", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"89", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"8f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"8f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"90", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"90", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"91", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"91", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"92", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"92", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"93", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"93", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"94", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"94", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"95", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"95", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"96", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"96", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"97", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"97", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"98", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"98", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"99", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"99", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9a", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9a", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9b", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9b", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9c", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9c", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9d", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9d", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9e", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9e", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"9f", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"9f", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"a9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"a9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"aa", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"aa", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ab", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ab", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ac", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ac", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ad", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ad", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ae", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ae", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"af", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"af", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"b9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"b9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ba", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ba", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"bb", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"bb", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"bc", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"bc", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"bd", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"bd", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"be", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"be", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"bf", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"bf", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"c9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"c9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ca", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ca", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"cb", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"cb", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"cc", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"cc", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"cd", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"cd", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ce", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ce", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"cf", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"cf", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"d9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"d9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"da", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"da", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"db", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"db", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"dc", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"dc", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"dd", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"dd", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"de", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"de", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"df", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"df", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"e9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"e9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ea", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ea", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"eb", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"eb", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ec", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ec", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ed", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ed", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ee", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ee", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ef", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ef", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f0", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f0", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f1", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f1", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f2", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f2", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f3", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f3", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f4", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f4", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f5", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f5", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f6", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f6", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f7", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f7", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f8", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f8", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"f9", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"f9", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"fa", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"fa", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"fb", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"fb", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"fc", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"fc", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"fd", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"fd", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"fe", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"fe", delay => 60),
    ( address => x"D0E2", write_p => '0', value => x"ff", delay => 2),
    ( address => x"D0E2", write_p => '1', value => x"ff", delay => 60),

    
    -- End of procedure
    others => ( address => x"FFFF", write_p => '0', value => x"00", delay => 1000)

    );

  signal idle_wait : integer := 0;
  
  signal expect_value : std_logic := '0';
  signal expected_value : unsigned(7 downto 0) := x"00";
  
begin

  buffered_uart0 : entity work.buffereduart port map (
    clock => cpuclock,
    reset => reset,
    irq => uart_irq,
    buffereduart_cs => buffereduart_cs,

    ---------------------------------------------------------------------------
    -- IO lines to the buffered UART
    ---------------------------------------------------------------------------
    uart_rx => buffereduart_rx,
    uart_tx => buffereduart_tx,
    uart_ringindicate => buffereduart_ringindicate,

    fastio_addr => unsigned(fastio_addr),
    fastio_write => fastio_write,
    fastio_read => fastio_read,
    fastio_rdata => fastio_rdata,
    fastio_wdata => fastio_wdata
    );

  
  process is
  begin
    -- pretend clock at 50MHz, just so the ns display is easier to read in simulation
    cpuclock <= '0';
    wait for 10 ns;
    cpuclock <= '1';
    wait for 10 ns;
  end process;
  
  
  process (cpuclock) is
  begin

    if rising_edge(cpuclock) then

      expect_value <= '0';
      fastio_read <= '0';
      fastio_write <= '0';
      
      if idle_wait /= 0 then
        idle_wait <= idle_wait - 1;
      else
        
        if mem_jobs(cycles).address = x"FFFF" then
          idle_wait <= mem_jobs(cycles).delay;
          expect_value <= '0';
          cycles <= 0;
          start_time <= current_time;          
        else
          cycles <= cycles + 1;        
          
          fastio_addr(15 downto 0) <= mem_jobs(cycles).address;
          fastio_addr(19 downto 16) <= x"0";
          fastio_read <= not mem_jobs(cycles).write_p;
          fastio_write <= mem_jobs(cycles).write_p;
          fastio_wdata <= mem_jobs(cycles).value;
          idle_wait <= mem_jobs(cycles).delay;
          
          if start_time = 0 then
            start_time <= current_time;
          end if;
          if (mem_jobs(cycles).write_p='0') then
            report "DISPATCHER: Reading from $" & to_hstring(mem_jobs(cycles).address) & ", expecting to see $"
              & to_hstring(mem_jobs(cycles).value);
            expect_value <= '1';
            expected_value <= mem_jobs(cycles).value;
          else
            report "DISPATCHER: Writing to $" & to_hstring(mem_jobs(cycles).address) & " <- $"
              & to_hstring(mem_jobs(cycles).value);
            expect_value <= '0';
            dispatch_time <= current_time;
          end if;
        end if;
      end if;
        
      if expect_value='1' then
        if fastio_rdata /= expected_value then
          report "DISPATCHER: ERROR: Read value $" & to_hstring(fastio_rdata) & ", expected to see $"
            & to_hstring(expected_value);
        else
          report "DISPATCHER: Read correct value $" & to_hstring(fastio_rdata);
        end if;
      end if;        
      
    end if;
      
  end process;
      
      
end foo;
     
