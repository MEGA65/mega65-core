library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-------------------------------------------------------------------------------

entity sid_tables is
	port (
          clock : in std_logic;
          sawtooth : in unsigned(11 downto 0);
          triangle : in unsigned(11 downto 0);
          st_out : out unsigned(7 downto 0) := x"00";
          p_t_out : out unsigned(7 downto 0) := x"00";
          ps_out : out unsigned(7 downto 0) := x"00";
          pst_out : out unsigned(7 downto 0) := x"00"
          );
end sid_tables;

architecture sequential of sid_tables is

begin

  process (clock,sawtooth,triangle) is
  begin
    if rising_edge(clock) then
      if sawtooth < x"07e" then   st_out <= x"00";
      elsif sawtooth < x"080" then   st_out <= x"03";
      elsif sawtooth < x"0fc" then   st_out <= x"00";
      elsif sawtooth < x"100" then   st_out <= x"07";
      elsif sawtooth < x"17e" then   st_out <= x"00";
      elsif sawtooth < x"180" then   st_out <= x"03";
      elsif sawtooth < x"1f8" then   st_out <= x"00";
      elsif sawtooth < x"1fc" then   st_out <= x"0e";
      elsif sawtooth < x"200" then   st_out <= x"0f";
      elsif sawtooth < x"27e" then   st_out <= x"00";
      elsif sawtooth < x"280" then   st_out <= x"03";
      elsif sawtooth < x"2fc" then   st_out <= x"00";
      elsif sawtooth < x"300" then   st_out <= x"07";
      elsif sawtooth < x"37e" then   st_out <= x"00";
      elsif sawtooth < x"380" then   st_out <= x"03";
      elsif sawtooth < x"3bf" then   st_out <= x"00";
      elsif sawtooth < x"3c0" then   st_out <= x"01";
      elsif sawtooth < x"3f0" then   st_out <= x"00";
      elsif sawtooth < x"3f8" then   st_out <= x"1c";
      elsif sawtooth < x"3fa" then   st_out <= x"1e";
      elsif sawtooth < x"400" then   st_out <= x"1f";
      elsif sawtooth < x"47e" then   st_out <= x"00";
      elsif sawtooth < x"480" then   st_out <= x"03";
      elsif sawtooth < x"4fc" then   st_out <= x"00";
      elsif sawtooth < x"500" then   st_out <= x"07";
      elsif sawtooth < x"57e" then   st_out <= x"00";
      elsif sawtooth < x"580" then   st_out <= x"03";
      elsif sawtooth < x"5f8" then   st_out <= x"00";
      elsif sawtooth < x"5fc" then   st_out <= x"0e";
      elsif sawtooth < x"5ff" then   st_out <= x"0f";
      elsif sawtooth < x"600" then   st_out <= x"1f";
      elsif sawtooth < x"67e" then   st_out <= x"00";
      elsif sawtooth < x"680" then   st_out <= x"03";
      elsif sawtooth < x"6fc" then   st_out <= x"00";
      elsif sawtooth < x"700" then   st_out <= x"07";
      elsif sawtooth < x"77e" then   st_out <= x"00";
      elsif sawtooth < x"780" then   st_out <= x"03";
      elsif sawtooth < x"7bf" then   st_out <= x"00";
      elsif sawtooth < x"7c0" then   st_out <= x"01";
      elsif sawtooth < x"7e0" then   st_out <= x"00";
      elsif sawtooth < x"7f0" then   st_out <= x"38";
      elsif sawtooth < x"7f7" then   st_out <= x"3c";
      elsif sawtooth < x"7f8" then   st_out <= x"3e";
      elsif sawtooth < x"800" then   st_out <= x"7f";
      elsif sawtooth < x"87e" then   st_out <= x"00";
      elsif sawtooth < x"880" then   st_out <= x"03";
      elsif sawtooth < x"8fc" then   st_out <= x"00";
      elsif sawtooth < x"900" then   st_out <= x"07";
      elsif sawtooth < x"97e" then   st_out <= x"00";
      elsif sawtooth < x"980" then   st_out <= x"03";
      elsif sawtooth < x"9f8" then   st_out <= x"00";
      elsif sawtooth < x"9fc" then   st_out <= x"0e";
      elsif sawtooth < x"a00" then   st_out <= x"0f";
      elsif sawtooth < x"a7e" then   st_out <= x"00";
      elsif sawtooth < x"a80" then   st_out <= x"03";
      elsif sawtooth < x"afc" then   st_out <= x"00";
      elsif sawtooth < x"b00" then   st_out <= x"07";
      elsif sawtooth < x"b7e" then   st_out <= x"00";
      elsif sawtooth < x"b80" then   st_out <= x"03";
      elsif sawtooth < x"bbf" then   st_out <= x"00";
      elsif sawtooth < x"bc0" then   st_out <= x"01";
      elsif sawtooth < x"bf0" then   st_out <= x"00";
      elsif sawtooth < x"bf8" then   st_out <= x"1c";
      elsif sawtooth < x"bfa" then   st_out <= x"1e";
      elsif sawtooth < x"bfe" then   st_out <= x"1f";
      elsif sawtooth < x"c00" then   st_out <= x"3f";
      elsif sawtooth < x"c7e" then   st_out <= x"00";
      elsif sawtooth < x"c80" then   st_out <= x"03";
      elsif sawtooth < x"cfc" then   st_out <= x"00";
      elsif sawtooth < x"d00" then   st_out <= x"07";
      elsif sawtooth < x"d7e" then   st_out <= x"00";
      elsif sawtooth < x"d80" then   st_out <= x"03";
      elsif sawtooth < x"dbf" then   st_out <= x"00";
      elsif sawtooth < x"dc0" then   st_out <= x"01";
      elsif sawtooth < x"df8" then   st_out <= x"00";
      elsif sawtooth < x"dfc" then   st_out <= x"0e";
      elsif sawtooth < x"dfe" then   st_out <= x"0f";
      elsif sawtooth < x"e00" then   st_out <= x"1f";
      elsif sawtooth < x"e7c" then   st_out <= x"00";
      elsif sawtooth < x"e7d" then   st_out <= x"80";
      elsif sawtooth < x"e7e" then   st_out <= x"00";
      elsif sawtooth < x"e80" then   st_out <= x"83";
      elsif sawtooth < x"efc" then   st_out <= x"80";
      elsif sawtooth < x"eff" then   st_out <= x"87";
      elsif sawtooth < x"f00" then   st_out <= x"8f";
      elsif sawtooth < x"f01" then   st_out <= x"c0";
      elsif sawtooth < x"f03" then   st_out <= x"e0";
      elsif sawtooth < x"f05" then   st_out <= x"c0";
      elsif sawtooth < x"f09" then   st_out <= x"e0";
      elsif sawtooth < x"f11" then   st_out <= x"c0";
      elsif sawtooth < x"f13" then   st_out <= x"e0";
      elsif sawtooth < x"f18" then   st_out <= x"c0";
      elsif sawtooth < x"f19" then   st_out <= x"e0";
      elsif sawtooth < x"f21" then   st_out <= x"c0";
      elsif sawtooth < x"f23" then   st_out <= x"e0";
      elsif sawtooth < x"f25" then   st_out <= x"c0";
      elsif sawtooth < x"f2b" then   st_out <= x"e0";
      elsif sawtooth < x"f2c" then   st_out <= x"c0";
      elsif sawtooth < x"f2d" then   st_out <= x"e0";
      elsif sawtooth < x"f2e" then   st_out <= x"c0";
      elsif sawtooth < x"f7e" then   st_out <= x"e0";
      elsif sawtooth < x"f80" then   st_out <= x"e3";
      elsif sawtooth < x"fbf" then   st_out <= x"f0";
      elsif sawtooth < x"fc0" then   st_out <= x"f1";
      elsif sawtooth < x"fe0" then   st_out <= x"f8";
      elsif sawtooth < x"ff0" then   st_out <= x"fc";
      elsif sawtooth < x"ff8" then   st_out <= x"fe";
      else  st_out <= x"ff";
      end if;

      if triangle(11 downto 1) < x"0ff" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"100" then   p_t_out <= x"07";
      elsif triangle(11 downto 1) < x"1fb" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"1fc" then   p_t_out <= x"1c";
      elsif triangle(11 downto 1) < x"1fd" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"1fe" then   p_t_out <= x"3c";
      elsif triangle(11 downto 1) < x"200" then   p_t_out <= x"3f";
      elsif triangle(11 downto 1) < x"2fd" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"2fe" then   p_t_out <= x"0c";
      elsif triangle(11 downto 1) < x"2ff" then   p_t_out <= x"5e";
      elsif triangle(11 downto 1) < x"300" then   p_t_out <= x"5f";
      elsif triangle(11 downto 1) < x"377" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"378" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"37b" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"37d" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"37f" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"380" then   p_t_out <= x"6f";
      elsif triangle(11 downto 1) < x"39f" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"3a0" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3ae" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"3b0" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3b3" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"3b7" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3b8" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3ba" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3be" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3bf" then   p_t_out <= x"70";
      elsif triangle(11 downto 1) < x"3c0" then   p_t_out <= x"77";
      elsif triangle(11 downto 1) < x"3c5" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"3cd" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3d0" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3d3" then   p_t_out <= x"40";
      elsif triangle(11 downto 1) < x"3d7" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3d8" then   p_t_out <= x"70";
      elsif triangle(11 downto 1) < x"3db" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3de" then   p_t_out <= x"70";
      elsif triangle(11 downto 1) < x"3df" then   p_t_out <= x"78";
      elsif triangle(11 downto 1) < x"3e0" then   p_t_out <= x"7b";
      elsif triangle(11 downto 1) < x"3e3" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3e4" then   p_t_out <= x"70";
      elsif triangle(11 downto 1) < x"3e5" then   p_t_out <= x"60";
      elsif triangle(11 downto 1) < x"3eb" then   p_t_out <= x"70";
      elsif triangle(11 downto 1) < x"3ef" then   p_t_out <= x"78";
      elsif triangle(11 downto 1) < x"3f0" then   p_t_out <= x"7c";
      elsif triangle(11 downto 1) < x"3f3" then   p_t_out <= x"78";
      elsif triangle(11 downto 1) < x"3f4" then   p_t_out <= x"7c";
      elsif triangle(11 downto 1) < x"3f5" then   p_t_out <= x"78";
      elsif triangle(11 downto 1) < x"3f7" then   p_t_out <= x"7c";
      elsif triangle(11 downto 1) < x"3f8" then   p_t_out <= x"7e";
      elsif triangle(11 downto 1) < x"3f9" then   p_t_out <= x"7c";
      elsif triangle(11 downto 1) < x"3fb" then   p_t_out <= x"7e";
      elsif triangle(11 downto 1) < x"400" then   p_t_out <= x"7f";
      elsif triangle(11 downto 1) < x"47f" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"480" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4bd" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"4c0" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4cf" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"4d0" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4d7" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"4d8" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4da" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"4e0" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4e3" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"4fe" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"4ff" then   p_t_out <= x"8e";
      elsif triangle(11 downto 1) < x"500" then   p_t_out <= x"9f";
      elsif triangle(11 downto 1) < x"51f" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"520" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"52b" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"52c" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"52d" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"530" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"532" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"540" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"543" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"544" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"545" then   p_t_out <= x"00";
      elsif triangle(11 downto 1) < x"57f" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"580" then   p_t_out <= x"af";
      elsif triangle(11 downto 1) < x"5bb" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"5bf" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5c0" then   p_t_out <= x"b7";
      elsif triangle(11 downto 1) < x"5cf" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"5d0" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5d6" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"5db" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5dc" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5dd" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5df" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5e0" then   p_t_out <= x"bb";
      elsif triangle(11 downto 1) < x"5e6" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5e8" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5e9" then   p_t_out <= x"a0";
      elsif triangle(11 downto 1) < x"5eb" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5ec" then   p_t_out <= x"b8";
      elsif triangle(11 downto 1) < x"5ed" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5ef" then   p_t_out <= x"b8";
      elsif triangle(11 downto 1) < x"5f0" then   p_t_out <= x"bc";
      elsif triangle(11 downto 1) < x"5f1" then   p_t_out <= x"b0";
      elsif triangle(11 downto 1) < x"5f5" then   p_t_out <= x"b8";
      elsif triangle(11 downto 1) < x"5f7" then   p_t_out <= x"bc";
      elsif triangle(11 downto 1) < x"5f8" then   p_t_out <= x"be";
      elsif triangle(11 downto 1) < x"5fa" then   p_t_out <= x"bc";
      elsif triangle(11 downto 1) < x"5fb" then   p_t_out <= x"be";
      elsif triangle(11 downto 1) < x"5fc" then   p_t_out <= x"bf";
      elsif triangle(11 downto 1) < x"5fd" then   p_t_out <= x"be";
      elsif triangle(11 downto 1) < x"600" then   p_t_out <= x"bf";
      elsif triangle(11 downto 1) < x"63e" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"640" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"657" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"658" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"65a" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"660" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"663" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"664" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"665" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"67f" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"680" then   p_t_out <= x"cf";
      elsif triangle(11 downto 1) < x"686" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"689" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"68a" then   p_t_out <= x"80";
      elsif triangle(11 downto 1) < x"6bf" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"6c0" then   p_t_out <= x"d7";
      elsif triangle(11 downto 1) < x"6dd" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"6df" then   p_t_out <= x"d0";
      elsif triangle(11 downto 1) < x"6e0" then   p_t_out <= x"d9";
      elsif triangle(11 downto 1) < x"6e7" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"6e8" then   p_t_out <= x"d0";
      elsif triangle(11 downto 1) < x"6e9" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"6ed" then   p_t_out <= x"d0";
      elsif triangle(11 downto 1) < x"6ef" then   p_t_out <= x"d8";
      elsif triangle(11 downto 1) < x"6f0" then   p_t_out <= x"dc";
      elsif triangle(11 downto 1) < x"6f2" then   p_t_out <= x"d0";
      elsif triangle(11 downto 1) < x"6f5" then   p_t_out <= x"d8";
      elsif triangle(11 downto 1) < x"6f7" then   p_t_out <= x"dc";
      elsif triangle(11 downto 1) < x"6f8" then   p_t_out <= x"de";
      elsif triangle(11 downto 1) < x"6fa" then   p_t_out <= x"dc";
      elsif triangle(11 downto 1) < x"6fb" then   p_t_out <= x"de";
      elsif triangle(11 downto 1) < x"6fc" then   p_t_out <= x"df";
      elsif triangle(11 downto 1) < x"6fd" then   p_t_out <= x"de";
      elsif triangle(11 downto 1) < x"700" then   p_t_out <= x"df";
      elsif triangle(11 downto 1) < x"71b" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"71c" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"71d" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"720" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"727" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"728" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"72a" then   p_t_out <= x"c0";
      elsif triangle(11 downto 1) < x"73f" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"740" then   p_t_out <= x"e7";
      elsif triangle(11 downto 1) < x"75f" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"760" then   p_t_out <= x"e8";
      elsif triangle(11 downto 1) < x"76e" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"76f" then   p_t_out <= x"e8";
      elsif triangle(11 downto 1) < x"770" then   p_t_out <= x"ec";
      elsif triangle(11 downto 1) < x"773" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"776" then   p_t_out <= x"e8";
      elsif triangle(11 downto 1) < x"777" then   p_t_out <= x"ec";
      elsif triangle(11 downto 1) < x"778" then   p_t_out <= x"ee";
      elsif triangle(11 downto 1) < x"77b" then   p_t_out <= x"ec";
      elsif triangle(11 downto 1) < x"77d" then   p_t_out <= x"ee";
      elsif triangle(11 downto 1) < x"780" then   p_t_out <= x"ef";
      elsif triangle(11 downto 1) < x"78d" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"790" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"792" then   p_t_out <= x"e0";
      elsif triangle(11 downto 1) < x"7af" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"7b0" then   p_t_out <= x"f4";
      elsif triangle(11 downto 1) < x"7b7" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"7b8" then   p_t_out <= x"f4";
      elsif triangle(11 downto 1) < x"7b9" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"7bb" then   p_t_out <= x"f4";
      elsif triangle(11 downto 1) < x"7bd" then   p_t_out <= x"f6";
      elsif triangle(11 downto 1) < x"7c0" then   p_t_out <= x"f7";
      elsif triangle(11 downto 1) < x"7c3" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"7c4" then   p_t_out <= x"f8";
      elsif triangle(11 downto 1) < x"7c5" then   p_t_out <= x"f0";
      elsif triangle(11 downto 1) < x"7db" then   p_t_out <= x"f8";
      elsif triangle(11 downto 1) < x"7dd" then   p_t_out <= x"fa";
      elsif triangle(11 downto 1) < x"7e0" then   p_t_out <= x"fb";
      elsif triangle(11 downto 1) < x"7e1" then   p_t_out <= x"f8";
      elsif triangle(11 downto 1) < x"7ed" then   p_t_out <= x"fc";
      elsif triangle(11 downto 1) < x"7f0" then   p_t_out <= x"fd";
      elsif triangle(11 downto 1) < x"7f8" then   p_t_out <= x"fe";
      else p_t_out <= x"ff";
      end if;

      if sawtooth < x"07f" then   ps_out <= x"00";
      elsif sawtooth < x"080" then   ps_out <= x"03";
      elsif sawtooth < x"0bf" then   ps_out <= x"00";
      elsif sawtooth < x"0c0" then   ps_out <= x"01";
      elsif sawtooth < x"0ff" then   ps_out <= x"00";
      elsif sawtooth < x"100" then   ps_out <= x"0f";
      elsif sawtooth < x"17f" then   ps_out <= x"00";
      elsif sawtooth < x"180" then   ps_out <= x"07";
      elsif sawtooth < x"1bf" then   ps_out <= x"00";
      elsif sawtooth < x"1c0" then   ps_out <= x"03";
      elsif sawtooth < x"1df" then   ps_out <= x"00";
      elsif sawtooth < x"1e0" then   ps_out <= x"01";
      elsif sawtooth < x"1fd" then   ps_out <= x"00";
      elsif sawtooth < x"1ff" then   ps_out <= x"07";
      elsif sawtooth < x"200" then   ps_out <= x"1f";
      elsif sawtooth < x"27f" then   ps_out <= x"00";
      elsif sawtooth < x"280" then   ps_out <= x"03";
      elsif sawtooth < x"2bf" then   ps_out <= x"00";
      elsif sawtooth < x"2c0" then   ps_out <= x"03";
      elsif sawtooth < x"2df" then   ps_out <= x"00";
      elsif sawtooth < x"2e0" then   ps_out <= x"01";
      elsif sawtooth < x"2fe" then   ps_out <= x"00";
      elsif sawtooth < x"2ff" then   ps_out <= x"01";
      elsif sawtooth < x"300" then   ps_out <= x"0f";
      elsif sawtooth < x"33f" then   ps_out <= x"00";
      elsif sawtooth < x"340" then   ps_out <= x"01";
      elsif sawtooth < x"37f" then   ps_out <= x"00";
      elsif sawtooth < x"380" then   ps_out <= x"17";
      elsif sawtooth < x"3bf" then   ps_out <= x"00";
      elsif sawtooth < x"3c0" then   ps_out <= x"3b";
      elsif sawtooth < x"3df" then   ps_out <= x"00";
      elsif sawtooth < x"3e0" then   ps_out <= x"3d";
      elsif sawtooth < x"3ef" then   ps_out <= x"00";
      elsif sawtooth < x"3f0" then   ps_out <= x"3e";
      elsif sawtooth < x"3f7" then   ps_out <= x"00";
      elsif sawtooth < x"3f8" then   ps_out <= x"3f";
      elsif sawtooth < x"3f9" then   ps_out <= x"00";
      elsif sawtooth < x"3fa" then   ps_out <= x"0c";
      elsif sawtooth < x"3fb" then   ps_out <= x"1c";
      elsif sawtooth < x"3fc" then   ps_out <= x"3f";
      elsif sawtooth < x"3fd" then   ps_out <= x"1e";
      elsif sawtooth < x"400" then   ps_out <= x"3f";
      elsif sawtooth < x"47f" then   ps_out <= x"00";
      elsif sawtooth < x"480" then   ps_out <= x"03";
      elsif sawtooth < x"4bf" then   ps_out <= x"00";
      elsif sawtooth < x"4c0" then   ps_out <= x"01";
      elsif sawtooth < x"4ff" then   ps_out <= x"00";
      elsif sawtooth < x"500" then   ps_out <= x"0f";
      elsif sawtooth < x"53f" then   ps_out <= x"00";
      elsif sawtooth < x"540" then   ps_out <= x"01";
      elsif sawtooth < x"57f" then   ps_out <= x"00";
      elsif sawtooth < x"580" then   ps_out <= x"07";
      elsif sawtooth < x"5bf" then   ps_out <= x"00";
      elsif sawtooth < x"5c0" then   ps_out <= x"0b";
      elsif sawtooth < x"5df" then   ps_out <= x"00";
      elsif sawtooth < x"5e0" then   ps_out <= x"0a";
      elsif sawtooth < x"5ef" then   ps_out <= x"00";
      elsif sawtooth < x"5f0" then   ps_out <= x"5e";
      elsif sawtooth < x"5f7" then   ps_out <= x"00";
      elsif sawtooth < x"5f8" then   ps_out <= x"5f";
      elsif sawtooth < x"5fb" then   ps_out <= x"00";
      elsif sawtooth < x"5fc" then   ps_out <= x"5f";
      elsif sawtooth < x"5fd" then   ps_out <= x"0c";
      elsif sawtooth < x"600" then   ps_out <= x"5f";
      elsif sawtooth < x"63f" then   ps_out <= x"00";
      elsif sawtooth < x"640" then   ps_out <= x"01";
      elsif sawtooth < x"67f" then   ps_out <= x"00";
      elsif sawtooth < x"680" then   ps_out <= x"47";
      elsif sawtooth < x"6bf" then   ps_out <= x"00";
      elsif sawtooth < x"6c0" then   ps_out <= x"43";
      elsif sawtooth < x"6df" then   ps_out <= x"00";
      elsif sawtooth < x"6e0" then   ps_out <= x"65";
      elsif sawtooth < x"6ef" then   ps_out <= x"00";
      elsif sawtooth < x"6f0" then   ps_out <= x"6e";
      elsif sawtooth < x"6f7" then   ps_out <= x"00";
      elsif sawtooth < x"6f8" then   ps_out <= x"6f";
      elsif sawtooth < x"6f9" then   ps_out <= x"00";
      elsif sawtooth < x"6fb" then   ps_out <= x"40";
      elsif sawtooth < x"6fc" then   ps_out <= x"6f";
      elsif sawtooth < x"6fd" then   ps_out <= x"40";
      elsif sawtooth < x"700" then   ps_out <= x"6f";
      elsif sawtooth < x"73f" then   ps_out <= x"00";
      elsif sawtooth < x"740" then   ps_out <= x"63";
      elsif sawtooth < x"75e" then   ps_out <= x"00";
      elsif sawtooth < x"75f" then   ps_out <= x"40";
      elsif sawtooth < x"760" then   ps_out <= x"61";
      elsif sawtooth < x"767" then   ps_out <= x"00";
      elsif sawtooth < x"768" then   ps_out <= x"40";
      elsif sawtooth < x"76b" then   ps_out <= x"00";
      elsif sawtooth < x"76c" then   ps_out <= x"40";
      elsif sawtooth < x"76d" then   ps_out <= x"00";
      elsif sawtooth < x"76f" then   ps_out <= x"40";
      elsif sawtooth < x"770" then   ps_out <= x"70";
      elsif sawtooth < x"772" then   ps_out <= x"00";
      elsif sawtooth < x"777" then   ps_out <= x"40";
      elsif sawtooth < x"778" then   ps_out <= x"70";
      elsif sawtooth < x"779" then   ps_out <= x"40";
      elsif sawtooth < x"77b" then   ps_out <= x"60";
      elsif sawtooth < x"77c" then   ps_out <= x"77";
      elsif sawtooth < x"77d" then   ps_out <= x"60";
      elsif sawtooth < x"780" then   ps_out <= x"77";
      elsif sawtooth < x"78f" then   ps_out <= x"00";
      elsif sawtooth < x"790" then   ps_out <= x"40";
      elsif sawtooth < x"796" then   ps_out <= x"00";
      elsif sawtooth < x"797" then   ps_out <= x"40";
      elsif sawtooth < x"798" then   ps_out <= x"60";
      elsif sawtooth < x"799" then   ps_out <= x"00";
      elsif sawtooth < x"79b" then   ps_out <= x"40";
      elsif sawtooth < x"79c" then   ps_out <= x"60";
      elsif sawtooth < x"79d" then   ps_out <= x"40";
      elsif sawtooth < x"79f" then   ps_out <= x"60";
      elsif sawtooth < x"7a0" then   ps_out <= x"79";
      elsif sawtooth < x"7a1" then   ps_out <= x"00";
      elsif sawtooth < x"7a7" then   ps_out <= x"40";
      elsif sawtooth < x"7a8" then   ps_out <= x"60";
      elsif sawtooth < x"7ab" then   ps_out <= x"40";
      elsif sawtooth < x"7af" then   ps_out <= x"60";
      elsif sawtooth < x"7b0" then   ps_out <= x"78";
      elsif sawtooth < x"7b1" then   ps_out <= x"40";
      elsif sawtooth < x"7b7" then   ps_out <= x"60";
      elsif sawtooth < x"7b8" then   ps_out <= x"78";
      elsif sawtooth < x"7b9" then   ps_out <= x"60";
      elsif sawtooth < x"7bb" then   ps_out <= x"70";
      elsif sawtooth < x"7bc" then   ps_out <= x"78";
      elsif sawtooth < x"7bd" then   ps_out <= x"70";
      elsif sawtooth < x"7be" then   ps_out <= x"79";
      elsif sawtooth < x"7c0" then   ps_out <= x"7b";
      elsif sawtooth < x"7c7" then   ps_out <= x"60";
      elsif sawtooth < x"7c8" then   ps_out <= x"70";
      elsif sawtooth < x"7cb" then   ps_out <= x"60";
      elsif sawtooth < x"7cc" then   ps_out <= x"70";
      elsif sawtooth < x"7cd" then   ps_out <= x"60";
      elsif sawtooth < x"7cf" then   ps_out <= x"70";
      elsif sawtooth < x"7d0" then   ps_out <= x"7c";
      elsif sawtooth < x"7d1" then   ps_out <= x"60";
      elsif sawtooth < x"7d7" then   ps_out <= x"70";
      elsif sawtooth < x"7d8" then   ps_out <= x"7c";
      elsif sawtooth < x"7d9" then   ps_out <= x"70";
      elsif sawtooth < x"7db" then   ps_out <= x"78";
      elsif sawtooth < x"7dc" then   ps_out <= x"7c";
      elsif sawtooth < x"7dd" then   ps_out <= x"78";
      elsif sawtooth < x"7df" then   ps_out <= x"7c";
      elsif sawtooth < x"7e0" then   ps_out <= x"7d";
      elsif sawtooth < x"7e1" then   ps_out <= x"70";
      elsif sawtooth < x"7e7" then   ps_out <= x"78";
      elsif sawtooth < x"7e8" then   ps_out <= x"7c";
      elsif sawtooth < x"7e9" then   ps_out <= x"78";
      elsif sawtooth < x"7eb" then   ps_out <= x"7c";
      elsif sawtooth < x"7ec" then   ps_out <= x"7e";
      elsif sawtooth < x"7ed" then   ps_out <= x"7c";
      elsif sawtooth < x"7f0" then   ps_out <= x"7e";
      elsif sawtooth < x"7f3" then   ps_out <= x"7c";
      elsif sawtooth < x"7f5" then   ps_out <= x"7e";
      elsif sawtooth < x"7f8" then   ps_out <= x"7f";
      elsif sawtooth < x"7f9" then   ps_out <= x"7e";
      elsif sawtooth < x"7ff" then   ps_out <= x"7f";
      elsif sawtooth < x"800" then   ps_out <= x"ff";
      elsif sawtooth < x"87f" then   ps_out <= x"00";
      elsif sawtooth < x"880" then   ps_out <= x"03";
      elsif sawtooth < x"8bf" then   ps_out <= x"00";
      elsif sawtooth < x"8c0" then   ps_out <= x"01";
      elsif sawtooth < x"8ff" then   ps_out <= x"00";
      elsif sawtooth < x"900" then   ps_out <= x"8f";
      elsif sawtooth < x"93f" then   ps_out <= x"00";
      elsif sawtooth < x"940" then   ps_out <= x"01";
      elsif sawtooth < x"97f" then   ps_out <= x"00";
      elsif sawtooth < x"980" then   ps_out <= x"87";
      elsif sawtooth < x"9bf" then   ps_out <= x"00";
      elsif sawtooth < x"9c0" then   ps_out <= x"83";
      elsif sawtooth < x"9de" then   ps_out <= x"00";
      elsif sawtooth < x"9df" then   ps_out <= x"80";
      elsif sawtooth < x"9e0" then   ps_out <= x"8d";
      elsif sawtooth < x"9e7" then   ps_out <= x"00";
      elsif sawtooth < x"9e8" then   ps_out <= x"80";
      elsif sawtooth < x"9eb" then   ps_out <= x"00";
      elsif sawtooth < x"9ec" then   ps_out <= x"80";
      elsif sawtooth < x"9ed" then   ps_out <= x"00";
      elsif sawtooth < x"9ef" then   ps_out <= x"80";
      elsif sawtooth < x"9f0" then   ps_out <= x"8e";
      elsif sawtooth < x"9f3" then   ps_out <= x"00";
      elsif sawtooth < x"9f7" then   ps_out <= x"80";
      elsif sawtooth < x"9f8" then   ps_out <= x"8f";
      elsif sawtooth < x"9fb" then   ps_out <= x"80";
      elsif sawtooth < x"9fc" then   ps_out <= x"9f";
      elsif sawtooth < x"9fd" then   ps_out <= x"80";
      elsif sawtooth < x"a00" then   ps_out <= x"9f";
      elsif sawtooth < x"a3f" then   ps_out <= x"00";
      elsif sawtooth < x"a40" then   ps_out <= x"01";
      elsif sawtooth < x"a6f" then   ps_out <= x"00";
      elsif sawtooth < x"a70" then   ps_out <= x"80";
      elsif sawtooth < x"a77" then   ps_out <= x"00";
      elsif sawtooth < x"a78" then   ps_out <= x"80";
      elsif sawtooth < x"a7b" then   ps_out <= x"00";
      elsif sawtooth < x"a7c" then   ps_out <= x"80";
      elsif sawtooth < x"a7d" then   ps_out <= x"00";
      elsif sawtooth < x"a7f" then   ps_out <= x"80";
      elsif sawtooth < x"a80" then   ps_out <= x"87";
      elsif sawtooth < x"a9f" then   ps_out <= x"00";
      elsif sawtooth < x"aa0" then   ps_out <= x"80";
      elsif sawtooth < x"aaf" then   ps_out <= x"00";
      elsif sawtooth < x"ab0" then   ps_out <= x"80";
      elsif sawtooth < x"ab7" then   ps_out <= x"00";
      elsif sawtooth < x"ab8" then   ps_out <= x"80";
      elsif sawtooth < x"abb" then   ps_out <= x"00";
      elsif sawtooth < x"abf" then   ps_out <= x"80";
      elsif sawtooth < x"ac0" then   ps_out <= x"83";
      elsif sawtooth < x"acf" then   ps_out <= x"00";
      elsif sawtooth < x"ad0" then   ps_out <= x"80";
      elsif sawtooth < x"ad5" then   ps_out <= x"00";
      elsif sawtooth < x"ad8" then   ps_out <= x"80";
      elsif sawtooth < x"ad9" then   ps_out <= x"00";
      elsif sawtooth < x"adf" then   ps_out <= x"80";
      elsif sawtooth < x"ae0" then   ps_out <= x"81";
      elsif sawtooth < x"aef" then   ps_out <= x"80";
      elsif sawtooth < x"af0" then   ps_out <= x"84";
      elsif sawtooth < x"af7" then   ps_out <= x"80";
      elsif sawtooth < x"af8" then   ps_out <= x"87";
      elsif sawtooth < x"afb" then   ps_out <= x"80";
      elsif sawtooth < x"afc" then   ps_out <= x"87";
      elsif sawtooth < x"afd" then   ps_out <= x"80";
      elsif sawtooth < x"afe" then   ps_out <= x"8f";
      elsif sawtooth < x"b00" then   ps_out <= x"af";
      elsif sawtooth < x"b0f" then   ps_out <= x"00";
      elsif sawtooth < x"b10" then   ps_out <= x"80";
      elsif sawtooth < x"b17" then   ps_out <= x"00";
      elsif sawtooth < x"b18" then   ps_out <= x"80";
      elsif sawtooth < x"b1b" then   ps_out <= x"00";
      elsif sawtooth < x"b20" then   ps_out <= x"80";
      elsif sawtooth < x"b23" then   ps_out <= x"00";
      elsif sawtooth < x"b24" then   ps_out <= x"80";
      elsif sawtooth < x"b26" then   ps_out <= x"00";
      elsif sawtooth < x"b28" then   ps_out <= x"80";
      elsif sawtooth < x"b29" then   ps_out <= x"00";
      elsif sawtooth < x"b3f" then   ps_out <= x"80";
      elsif sawtooth < x"b40" then   ps_out <= x"83";
      elsif sawtooth < x"b5f" then   ps_out <= x"80";
      elsif sawtooth < x"b60" then   ps_out <= x"81";
      elsif sawtooth < x"b6f" then   ps_out <= x"80";
      elsif sawtooth < x"b70" then   ps_out <= x"a0";
      elsif sawtooth < x"b77" then   ps_out <= x"80";
      elsif sawtooth < x"b78" then   ps_out <= x"a0";
      elsif sawtooth < x"b7b" then   ps_out <= x"80";
      elsif sawtooth < x"b7c" then   ps_out <= x"a0";
      elsif sawtooth < x"b7d" then   ps_out <= x"80";
      elsif sawtooth < x"b7e" then   ps_out <= x"a3";
      elsif sawtooth < x"b80" then   ps_out <= x"b7";
      elsif sawtooth < x"b9f" then   ps_out <= x"80";
      elsif sawtooth < x"ba0" then   ps_out <= x"b1";
      elsif sawtooth < x"baf" then   ps_out <= x"80";
      elsif sawtooth < x"bb0" then   ps_out <= x"b0";
      elsif sawtooth < x"bb7" then   ps_out <= x"80";
      elsif sawtooth < x"bb8" then   ps_out <= x"b0";
      elsif sawtooth < x"bb9" then   ps_out <= x"80";
      elsif sawtooth < x"bbb" then   ps_out <= x"a0";
      elsif sawtooth < x"bbc" then   ps_out <= x"b0";
      elsif sawtooth < x"bbd" then   ps_out <= x"a0";
      elsif sawtooth < x"bbe" then   ps_out <= x"b8";
      elsif sawtooth < x"bbf" then   ps_out <= x"b9";
      elsif sawtooth < x"bc0" then   ps_out <= x"bb";
      elsif sawtooth < x"bc7" then   ps_out <= x"80";
      elsif sawtooth < x"bc8" then   ps_out <= x"a0";
      elsif sawtooth < x"bcb" then   ps_out <= x"80";
      elsif sawtooth < x"bcc" then   ps_out <= x"a0";
      elsif sawtooth < x"bcd" then   ps_out <= x"80";
      elsif sawtooth < x"bcf" then   ps_out <= x"a0";
      elsif sawtooth < x"bd0" then   ps_out <= x"b8";
      elsif sawtooth < x"bd1" then   ps_out <= x"80";
      elsif sawtooth < x"bd7" then   ps_out <= x"a0";
      elsif sawtooth < x"bd8" then   ps_out <= x"b8";
      elsif sawtooth < x"bd9" then   ps_out <= x"a0";
      elsif sawtooth < x"bdb" then   ps_out <= x"b0";
      elsif sawtooth < x"bdc" then   ps_out <= x"b8";
      elsif sawtooth < x"bdd" then   ps_out <= x"b0";
      elsif sawtooth < x"bdf" then   ps_out <= x"bc";
      elsif sawtooth < x"be0" then   ps_out <= x"bd";
      elsif sawtooth < x"be1" then   ps_out <= x"a0";
      elsif sawtooth < x"be5" then   ps_out <= x"b0";
      elsif sawtooth < x"be7" then   ps_out <= x"b8";
      elsif sawtooth < x"be8" then   ps_out <= x"bc";
      elsif sawtooth < x"be9" then   ps_out <= x"b0";
      elsif sawtooth < x"beb" then   ps_out <= x"b8";
      elsif sawtooth < x"bec" then   ps_out <= x"bc";
      elsif sawtooth < x"bed" then   ps_out <= x"b8";
      elsif sawtooth < x"bee" then   ps_out <= x"bc";
      elsif sawtooth < x"bf0" then   ps_out <= x"be";
      elsif sawtooth < x"bf1" then   ps_out <= x"b8";
      elsif sawtooth < x"bf3" then   ps_out <= x"bc";
      elsif sawtooth < x"bf4" then   ps_out <= x"be";
      elsif sawtooth < x"bf5" then   ps_out <= x"bc";
      elsif sawtooth < x"bf7" then   ps_out <= x"be";
      elsif sawtooth < x"bf8" then   ps_out <= x"bf";
      elsif sawtooth < x"bf9" then   ps_out <= x"be";
      elsif sawtooth < x"c00" then   ps_out <= x"bf";
      elsif sawtooth < x"c03" then   ps_out <= x"00";
      elsif sawtooth < x"c04" then   ps_out <= x"80";
      elsif sawtooth < x"c07" then   ps_out <= x"00";
      elsif sawtooth < x"c08" then   ps_out <= x"80";
      elsif sawtooth < x"c0b" then   ps_out <= x"00";
      elsif sawtooth < x"c0c" then   ps_out <= x"80";
      elsif sawtooth < x"c0f" then   ps_out <= x"00";
      elsif sawtooth < x"c10" then   ps_out <= x"80";
      elsif sawtooth < x"c11" then   ps_out <= x"00";
      elsif sawtooth < x"c18" then   ps_out <= x"80";
      elsif sawtooth < x"c19" then   ps_out <= x"00";
      elsif sawtooth < x"c3f" then   ps_out <= x"80";
      elsif sawtooth < x"c40" then   ps_out <= x"81";
      elsif sawtooth < x"c7f" then   ps_out <= x"80";
      elsif sawtooth < x"c80" then   ps_out <= x"c7";
      elsif sawtooth < x"cbe" then   ps_out <= x"80";
      elsif sawtooth < x"cbf" then   ps_out <= x"c0";
      elsif sawtooth < x"cc0" then   ps_out <= x"c3";
      elsif sawtooth < x"ccf" then   ps_out <= x"80";
      elsif sawtooth < x"cd0" then   ps_out <= x"c0";
      elsif sawtooth < x"cd7" then   ps_out <= x"80";
      elsif sawtooth < x"cd8" then   ps_out <= x"c0";
      elsif sawtooth < x"cdb" then   ps_out <= x"80";
      elsif sawtooth < x"cdc" then   ps_out <= x"c0";
      elsif sawtooth < x"cdd" then   ps_out <= x"80";
      elsif sawtooth < x"cdf" then   ps_out <= x"c0";
      elsif sawtooth < x"ce0" then   ps_out <= x"c1";
      elsif sawtooth < x"ce7" then   ps_out <= x"80";
      elsif sawtooth < x"ce8" then   ps_out <= x"c0";
      elsif sawtooth < x"ceb" then   ps_out <= x"80";
      elsif sawtooth < x"cf7" then   ps_out <= x"c0";
      elsif sawtooth < x"cf8" then   ps_out <= x"c7";
      elsif sawtooth < x"cfb" then   ps_out <= x"c0";
      elsif sawtooth < x"cfc" then   ps_out <= x"c7";
      elsif sawtooth < x"cfd" then   ps_out <= x"c0";
      elsif sawtooth < x"d00" then   ps_out <= x"cf";
      elsif sawtooth < x"d1f" then   ps_out <= x"80";
      elsif sawtooth < x"d20" then   ps_out <= x"c0";
      elsif sawtooth < x"d2f" then   ps_out <= x"80";
      elsif sawtooth < x"d30" then   ps_out <= x"c0";
      elsif sawtooth < x"d36" then   ps_out <= x"80";
      elsif sawtooth < x"d38" then   ps_out <= x"c0";
      elsif sawtooth < x"d39" then   ps_out <= x"80";
      elsif sawtooth < x"d3f" then   ps_out <= x"c0";
      elsif sawtooth < x"d40" then   ps_out <= x"c3";
      elsif sawtooth < x"d47" then   ps_out <= x"80";
      elsif sawtooth < x"d48" then   ps_out <= x"c0";
      elsif sawtooth < x"d4b" then   ps_out <= x"80";
      elsif sawtooth < x"d4c" then   ps_out <= x"c0";
      elsif sawtooth < x"d4d" then   ps_out <= x"80";
      elsif sawtooth < x"d50" then   ps_out <= x"c0";
      elsif sawtooth < x"d51" then   ps_out <= x"80";
      elsif sawtooth < x"d5f" then   ps_out <= x"c0";
      elsif sawtooth < x"d60" then   ps_out <= x"c1";
      elsif sawtooth < x"d7d" then   ps_out <= x"c0";
      elsif sawtooth < x"d7e" then   ps_out <= x"c1";
      elsif sawtooth < x"d7f" then   ps_out <= x"c7";
      elsif sawtooth < x"d80" then   ps_out <= x"d7";
      elsif sawtooth < x"daf" then   ps_out <= x"c0";
      elsif sawtooth < x"db0" then   ps_out <= x"d0";
      elsif sawtooth < x"db7" then   ps_out <= x"c0";
      elsif sawtooth < x"db8" then   ps_out <= x"d0";
      elsif sawtooth < x"dbb" then   ps_out <= x"c0";
      elsif sawtooth < x"dbc" then   ps_out <= x"d0";
      elsif sawtooth < x"dbd" then   ps_out <= x"c0";
      elsif sawtooth < x"dbe" then   ps_out <= x"d0";
      elsif sawtooth < x"dbf" then   ps_out <= x"d8";
      elsif sawtooth < x"dc0" then   ps_out <= x"db";
      elsif sawtooth < x"dcf" then   ps_out <= x"c0";
      elsif sawtooth < x"dd0" then   ps_out <= x"d8";
      elsif sawtooth < x"dd7" then   ps_out <= x"c0";
      elsif sawtooth < x"dd8" then   ps_out <= x"d8";
      elsif sawtooth < x"ddb" then   ps_out <= x"c0";
      elsif sawtooth < x"ddc" then   ps_out <= x"d8";
      elsif sawtooth < x"ddd" then   ps_out <= x"d0";
      elsif sawtooth < x"ddf" then   ps_out <= x"d8";
      elsif sawtooth < x"de0" then   ps_out <= x"dd";
      elsif sawtooth < x"de3" then   ps_out <= x"c0";
      elsif sawtooth < x"de4" then   ps_out <= x"d0";
      elsif sawtooth < x"de5" then   ps_out <= x"c0";
      elsif sawtooth < x"de7" then   ps_out <= x"d0";
      elsif sawtooth < x"de8" then   ps_out <= x"dc";
      elsif sawtooth < x"de9" then   ps_out <= x"d0";
      elsif sawtooth < x"deb" then   ps_out <= x"d8";
      elsif sawtooth < x"dec" then   ps_out <= x"dc";
      elsif sawtooth < x"ded" then   ps_out <= x"d8";
      elsif sawtooth < x"def" then   ps_out <= x"dc";
      elsif sawtooth < x"df0" then   ps_out <= x"de";
      elsif sawtooth < x"df1" then   ps_out <= x"d8";
      elsif sawtooth < x"df3" then   ps_out <= x"dc";
      elsif sawtooth < x"df4" then   ps_out <= x"de";
      elsif sawtooth < x"df5" then   ps_out <= x"dc";
      elsif sawtooth < x"df7" then   ps_out <= x"de";
      elsif sawtooth < x"df8" then   ps_out <= x"df";
      elsif sawtooth < x"df9" then   ps_out <= x"de";
      elsif sawtooth < x"e00" then   ps_out <= x"df";
      elsif sawtooth < x"e3f" then   ps_out <= x"c0";
      elsif sawtooth < x"e40" then   ps_out <= x"e3";
      elsif sawtooth < x"e57" then   ps_out <= x"c0";
      elsif sawtooth < x"e58" then   ps_out <= x"e0";
      elsif sawtooth < x"e5b" then   ps_out <= x"c0";
      elsif sawtooth < x"e5c" then   ps_out <= x"e0";
      elsif sawtooth < x"e5d" then   ps_out <= x"c0";
      elsif sawtooth < x"e5f" then   ps_out <= x"e0";
      elsif sawtooth < x"e60" then   ps_out <= x"e1";
      elsif sawtooth < x"e67" then   ps_out <= x"c0";
      elsif sawtooth < x"e68" then   ps_out <= x"e0";
      elsif sawtooth < x"e6b" then   ps_out <= x"c0";
      elsif sawtooth < x"e70" then   ps_out <= x"e0";
      elsif sawtooth < x"e71" then   ps_out <= x"c0";
      elsif sawtooth < x"e7d" then   ps_out <= x"e0";
      elsif sawtooth < x"e7e" then   ps_out <= x"e1";
      elsif sawtooth < x"e7f" then   ps_out <= x"e3";
      elsif sawtooth < x"e80" then   ps_out <= x"e7";
      elsif sawtooth < x"e87" then   ps_out <= x"c0";
      elsif sawtooth < x"e88" then   ps_out <= x"e0";
      elsif sawtooth < x"e8b" then   ps_out <= x"c0";
      elsif sawtooth < x"e8c" then   ps_out <= x"e0";
      elsif sawtooth < x"e8d" then   ps_out <= x"c0";
      elsif sawtooth < x"e90" then   ps_out <= x"e0";
      elsif sawtooth < x"e93" then   ps_out <= x"c0";
      elsif sawtooth < x"e94" then   ps_out <= x"e0";
      elsif sawtooth < x"e95" then   ps_out <= x"c0";
      elsif sawtooth < x"ebf" then   ps_out <= x"e0";
      elsif sawtooth < x"ec0" then   ps_out <= x"eb";
      elsif sawtooth < x"edb" then   ps_out <= x"e0";
      elsif sawtooth < x"edc" then   ps_out <= x"e8";
      elsif sawtooth < x"edd" then   ps_out <= x"e0";
      elsif sawtooth < x"edf" then   ps_out <= x"e8";
      elsif sawtooth < x"ee0" then   ps_out <= x"ed";
      elsif sawtooth < x"ee7" then   ps_out <= x"e0";
      elsif sawtooth < x"ee8" then   ps_out <= x"ec";
      elsif sawtooth < x"eeb" then   ps_out <= x"e0";
      elsif sawtooth < x"eec" then   ps_out <= x"ec";
      elsif sawtooth < x"eed" then   ps_out <= x"e8";
      elsif sawtooth < x"eef" then   ps_out <= x"ec";
      elsif sawtooth < x"ef0" then   ps_out <= x"ee";
      elsif sawtooth < x"ef3" then   ps_out <= x"e8";
      elsif sawtooth < x"ef5" then   ps_out <= x"ec";
      elsif sawtooth < x"ef7" then   ps_out <= x"ee";
      elsif sawtooth < x"ef8" then   ps_out <= x"ef";
      elsif sawtooth < x"ef9" then   ps_out <= x"ec";
      elsif sawtooth < x"f00" then   ps_out <= x"ef";
      elsif sawtooth < x"f1f" then   ps_out <= x"e0";
      elsif sawtooth < x"f20" then   ps_out <= x"f0";
      elsif sawtooth < x"f27" then   ps_out <= x"e0";
      elsif sawtooth < x"f28" then   ps_out <= x"f0";
      elsif sawtooth < x"f2b" then   ps_out <= x"e0";
      elsif sawtooth < x"f2c" then   ps_out <= x"f0";
      elsif sawtooth < x"f2d" then   ps_out <= x"e0";
      elsif sawtooth < x"f30" then   ps_out <= x"f0";
      elsif sawtooth < x"f33" then   ps_out <= x"e0";
      elsif sawtooth < x"f3f" then   ps_out <= x"f0";
      elsif sawtooth < x"f40" then   ps_out <= x"f3";
      elsif sawtooth < x"f43" then   ps_out <= x"e0";
      elsif sawtooth < x"f5f" then   ps_out <= x"f0";
      elsif sawtooth < x"f60" then   ps_out <= x"f5";
      elsif sawtooth < x"f6d" then   ps_out <= x"f0";
      elsif sawtooth < x"f6f" then   ps_out <= x"f4";
      elsif sawtooth < x"f70" then   ps_out <= x"f6";
      elsif sawtooth < x"f73" then   ps_out <= x"f0";
      elsif sawtooth < x"f74" then   ps_out <= x"f4";
      elsif sawtooth < x"f75" then   ps_out <= x"f0";
      elsif sawtooth < x"f76" then   ps_out <= x"f4";
      elsif sawtooth < x"f77" then   ps_out <= x"f6";
      elsif sawtooth < x"f78" then   ps_out <= x"f7";
      elsif sawtooth < x"f79" then   ps_out <= x"f4";
      elsif sawtooth < x"f7b" then   ps_out <= x"f6";
      elsif sawtooth < x"f80" then   ps_out <= x"f7";
      elsif sawtooth < x"f87" then   ps_out <= x"f0";
      elsif sawtooth < x"f88" then   ps_out <= x"f8";
      elsif sawtooth < x"f8d" then   ps_out <= x"f0";
      elsif sawtooth < x"f90" then   ps_out <= x"f8";
      elsif sawtooth < x"f93" then   ps_out <= x"f0";
      elsif sawtooth < x"f94" then   ps_out <= x"f8";
      elsif sawtooth < x"f95" then   ps_out <= x"f0";
      elsif sawtooth < x"f9f" then   ps_out <= x"f8";
      elsif sawtooth < x"fa0" then   ps_out <= x"f9";
      elsif sawtooth < x"faf" then   ps_out <= x"f8";
      elsif sawtooth < x"fb0" then   ps_out <= x"fa";
      elsif sawtooth < x"fb7" then   ps_out <= x"f8";
      elsif sawtooth < x"fb8" then   ps_out <= x"fb";
      elsif sawtooth < x"fb9" then   ps_out <= x"f8";
      elsif sawtooth < x"fbb" then   ps_out <= x"fa";
      elsif sawtooth < x"fc0" then   ps_out <= x"fb";
      elsif sawtooth < x"fc3" then   ps_out <= x"f8";
      elsif sawtooth < x"fc4" then   ps_out <= x"fc";
      elsif sawtooth < x"fc5" then   ps_out <= x"f8";
      elsif sawtooth < x"fd7" then   ps_out <= x"fc";
      elsif sawtooth < x"fd8" then   ps_out <= x"fd";
      elsif sawtooth < x"fdb" then   ps_out <= x"fc";
      elsif sawtooth < x"fe0" then   ps_out <= x"fd";
      elsif sawtooth < x"fe2" then   ps_out <= x"fc";
      elsif sawtooth < x"ff0" then   ps_out <= x"fe";
      else  ps_out <= x"ff";
      end if;

      if sawtooth < x"3ff" then   pst_out <= x"00";
      elsif sawtooth < x"400" then   pst_out <= x"1f";
      elsif sawtooth < x"7ee" then   pst_out <= x"00";
      elsif sawtooth < x"7ef" then   pst_out <= x"20";
      elsif sawtooth < x"7f0" then   pst_out <= x"70";
      elsif sawtooth < x"7f1" then   pst_out <= x"60";
      elsif sawtooth < x"7f2" then   pst_out <= x"20";
      elsif sawtooth < x"7f7" then   pst_out <= x"70";
      elsif sawtooth < x"7fa" then   pst_out <= x"78";
      elsif sawtooth < x"7fc" then   pst_out <= x"7c";
      elsif sawtooth < x"7fe" then   pst_out <= x"7e";
      elsif sawtooth < x"800" then   pst_out <= x"7f";
      elsif sawtooth < x"bfd" then   pst_out <= x"00";
      elsif sawtooth < x"bfe" then   pst_out <= x"08";
      elsif sawtooth < x"bff" then   pst_out <= x"1e";
      elsif sawtooth < x"c00" then   pst_out <= x"3f";
      elsif sawtooth < x"df7" then   pst_out <= x"00";
      elsif sawtooth < x"dfe" then   pst_out <= x"80";
      elsif sawtooth < x"dff" then   pst_out <= x"8c";
      elsif sawtooth < x"e00" then   pst_out <= x"9f";
      elsif sawtooth < x"e3e" then   pst_out <= x"00";
      elsif sawtooth < x"e40" then   pst_out <= x"80";
      elsif sawtooth < x"e5e" then   pst_out <= x"00";
      elsif sawtooth < x"e60" then   pst_out <= x"80";
      elsif sawtooth < x"e66" then   pst_out <= x"00";
      elsif sawtooth < x"e67" then   pst_out <= x"80";
      elsif sawtooth < x"e6a" then   pst_out <= x"00";
      elsif sawtooth < x"e80" then   pst_out <= x"80";
      elsif sawtooth < x"e82" then   pst_out <= x"00";
      elsif sawtooth < x"e83" then   pst_out <= x"80";
      elsif sawtooth < x"e85" then   pst_out <= x"00";
      elsif sawtooth < x"e89" then   pst_out <= x"80";
      elsif sawtooth < x"e8a" then   pst_out <= x"00";
      elsif sawtooth < x"eee" then   pst_out <= x"80";
      elsif sawtooth < x"eff" then   pst_out <= x"c0";
      elsif sawtooth < x"f00" then   pst_out <= x"cf";
      elsif sawtooth < x"f6f" then   pst_out <= x"c0";
      elsif sawtooth < x"f70" then   pst_out <= x"e0";
      elsif sawtooth < x"f74" then   pst_out <= x"c0";
      elsif sawtooth < x"f7f" then   pst_out <= x"e0";
      elsif sawtooth < x"f80" then   pst_out <= x"e3";
      elsif sawtooth < x"fb6" then   pst_out <= x"e0";
      elsif sawtooth < x"fda" then   pst_out <= x"f0";
      elsif sawtooth < x"feb" then   pst_out <= x"f8";
      elsif sawtooth < x"ff5" then   pst_out <= x"fc";
      elsif sawtooth < x"ff9" then   pst_out <= x"fe";
      else  pst_out <= x"ff";
      end if;
      
      
    end if;
  end process;
  
end sequential;
